
module SNPS_CLOCK_GATE_HIGH_input_fifo_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  TLATNTSCAX2 latch ( .E(EN), .SE(TE), .CK(CLK), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_input_fifo_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  TLATNTSCAX2 latch ( .E(EN), .SE(TE), .CK(CLK), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_input_fifo_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  TLATNTSCAX2 latch ( .E(EN), .SE(TE), .CK(CLK), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_input_fifo_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  TLATNTSCAX2 latch ( .E(EN), .SE(TE), .CK(CLK), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_input_fifo_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  TLATNTSCAX2 latch ( .E(EN), .SE(TE), .CK(CLK), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_input_fifo_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  TLATNTSCAX2 latch ( .E(EN), .SE(TE), .CK(CLK), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_input_fifo_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  TLATNTSCAX2 latch ( .E(EN), .SE(TE), .CK(CLK), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_input_fifo_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  TLATNTSCAX2 latch ( .E(EN), .SE(TE), .CK(CLK), .ECK(ENCLK) );
endmodule


module chip ( clk_PAD, rst_PAD, data_recv_PAD, data_dec_PAD );
  input [15:0] data_recv_PAD;
  output [7:0] data_dec_PAD;
  input clk_PAD, rst_PAD;
  wire   io_clk, io_rst, \decoder/w_PM_4[6] , \decoder/w_PM_3[6] ,
         \decoder/w_PM_2[6] , \decoder/w_PM_2[5] , \decoder/w_PM_1[6] ,
         \decoder/w_PM_1[5] , \decoder/w_PM_1[3] , \decoder/w_PM_1[1] ,
         \decoder/w_PM_1[0] , \decoder/w_data_4[6] , \decoder/w_data_4[5] ,
         \decoder/w_data_4[4] , \decoder/w_data_3[7] , \decoder/w_data_3[6] ,
         \decoder/w_data_3[5] , \decoder/w_data_3[4] , \decoder/w_data_3[3] ,
         \decoder/w_data_3[2] , \decoder/w_data_2[2] , \decoder/w_data_1[2] ,
         \decoder/w_enc_bit_8[0] , \decoder/w_enc_bit_7[0] ,
         \decoder/w_enc_bit_6[0] , \decoder/w_enc_bit_5[0] ,
         \decoder/w_enc_bit_4[0] , \decoder/w_enc_bit_3[0] ,
         \decoder/w_enc_bit_2[0] , \decoder/u_input_shifter/w_data_8[15] ,
         \decoder/u_input_shifter/w_data_8[14] ,
         \decoder/u_input_shifter/w_data_8[13] ,
         \decoder/u_input_shifter/w_data_8[12] ,
         \decoder/u_input_shifter/w_data_8[11] ,
         \decoder/u_input_shifter/w_data_8[10] ,
         \decoder/u_input_shifter/w_data_8[9] ,
         \decoder/u_input_shifter/w_data_8[8] ,
         \decoder/u_input_shifter/w_data_8[7] ,
         \decoder/u_input_shifter/w_data_8[6] ,
         \decoder/u_input_shifter/w_data_8[5] ,
         \decoder/u_input_shifter/w_data_8[4] ,
         \decoder/u_input_shifter/w_data_8[3] ,
         \decoder/u_input_shifter/w_data_8[2] ,
         \decoder/u_input_shifter/w_data_8[1] ,
         \decoder/u_input_shifter/w_data_8[0] ,
         \decoder/u_input_shifter/w_data_7[15] ,
         \decoder/u_input_shifter/w_data_7[14] ,
         \decoder/u_input_shifter/w_data_7[13] ,
         \decoder/u_input_shifter/w_data_7[12] ,
         \decoder/u_input_shifter/w_data_7[11] ,
         \decoder/u_input_shifter/w_data_7[10] ,
         \decoder/u_input_shifter/w_data_7[9] ,
         \decoder/u_input_shifter/w_data_7[8] ,
         \decoder/u_input_shifter/w_data_7[7] ,
         \decoder/u_input_shifter/w_data_7[6] ,
         \decoder/u_input_shifter/w_data_7[5] ,
         \decoder/u_input_shifter/w_data_7[4] ,
         \decoder/u_input_shifter/w_data_7[3] ,
         \decoder/u_input_shifter/w_data_7[2] ,
         \decoder/u_input_shifter/w_data_7[1] ,
         \decoder/u_input_shifter/w_data_7[0] ,
         \decoder/u_input_shifter/w_data_6[15] ,
         \decoder/u_input_shifter/w_data_6[14] ,
         \decoder/u_input_shifter/w_data_6[13] ,
         \decoder/u_input_shifter/w_data_6[12] ,
         \decoder/u_input_shifter/w_data_6[11] ,
         \decoder/u_input_shifter/w_data_6[10] ,
         \decoder/u_input_shifter/w_data_6[9] ,
         \decoder/u_input_shifter/w_data_6[8] ,
         \decoder/u_input_shifter/w_data_6[7] ,
         \decoder/u_input_shifter/w_data_6[6] ,
         \decoder/u_input_shifter/w_data_6[5] ,
         \decoder/u_input_shifter/w_data_6[4] ,
         \decoder/u_input_shifter/w_data_6[3] ,
         \decoder/u_input_shifter/w_data_6[2] ,
         \decoder/u_input_shifter/w_data_6[1] ,
         \decoder/u_input_shifter/w_data_6[0] ,
         \decoder/u_input_shifter/w_data_5[15] ,
         \decoder/u_input_shifter/w_data_5[14] ,
         \decoder/u_input_shifter/w_data_5[13] ,
         \decoder/u_input_shifter/w_data_5[12] ,
         \decoder/u_input_shifter/w_data_5[11] ,
         \decoder/u_input_shifter/w_data_5[10] ,
         \decoder/u_input_shifter/w_data_5[9] ,
         \decoder/u_input_shifter/w_data_5[8] ,
         \decoder/u_input_shifter/w_data_5[7] ,
         \decoder/u_input_shifter/w_data_5[6] ,
         \decoder/u_input_shifter/w_data_5[5] ,
         \decoder/u_input_shifter/w_data_5[4] ,
         \decoder/u_input_shifter/w_data_5[3] ,
         \decoder/u_input_shifter/w_data_5[2] ,
         \decoder/u_input_shifter/w_data_5[1] ,
         \decoder/u_input_shifter/w_data_5[0] ,
         \decoder/u_input_shifter/w_data_4[15] ,
         \decoder/u_input_shifter/w_data_4[14] ,
         \decoder/u_input_shifter/w_data_4[13] ,
         \decoder/u_input_shifter/w_data_4[12] ,
         \decoder/u_input_shifter/w_data_4[11] ,
         \decoder/u_input_shifter/w_data_4[10] ,
         \decoder/u_input_shifter/w_data_4[9] ,
         \decoder/u_input_shifter/w_data_4[8] ,
         \decoder/u_input_shifter/w_data_4[7] ,
         \decoder/u_input_shifter/w_data_4[6] ,
         \decoder/u_input_shifter/w_data_4[5] ,
         \decoder/u_input_shifter/w_data_4[4] ,
         \decoder/u_input_shifter/w_data_4[3] ,
         \decoder/u_input_shifter/w_data_4[2] ,
         \decoder/u_input_shifter/w_data_4[1] ,
         \decoder/u_input_shifter/w_data_4[0] ,
         \decoder/u_input_shifter/w_data_3[15] ,
         \decoder/u_input_shifter/w_data_3[14] ,
         \decoder/u_input_shifter/w_data_3[13] ,
         \decoder/u_input_shifter/w_data_3[12] ,
         \decoder/u_input_shifter/w_data_3[11] ,
         \decoder/u_input_shifter/w_data_3[10] ,
         \decoder/u_input_shifter/w_data_3[9] ,
         \decoder/u_input_shifter/w_data_3[8] ,
         \decoder/u_input_shifter/w_data_3[7] ,
         \decoder/u_input_shifter/w_data_3[6] ,
         \decoder/u_input_shifter/w_data_3[5] ,
         \decoder/u_input_shifter/w_data_3[4] ,
         \decoder/u_input_shifter/w_data_3[3] ,
         \decoder/u_input_shifter/w_data_3[2] ,
         \decoder/u_input_shifter/w_data_3[1] ,
         \decoder/u_input_shifter/w_data_3[0] ,
         \decoder/u_input_shifter/w_data_2[15] ,
         \decoder/u_input_shifter/w_data_2[14] ,
         \decoder/u_input_shifter/w_data_2[13] ,
         \decoder/u_input_shifter/w_data_2[12] ,
         \decoder/u_input_shifter/w_data_2[11] ,
         \decoder/u_input_shifter/w_data_2[10] ,
         \decoder/u_input_shifter/w_data_2[9] ,
         \decoder/u_input_shifter/w_data_2[8] ,
         \decoder/u_input_shifter/w_data_2[7] ,
         \decoder/u_input_shifter/w_data_2[6] ,
         \decoder/u_input_shifter/w_data_2[5] ,
         \decoder/u_input_shifter/w_data_2[4] ,
         \decoder/u_input_shifter/w_data_2[3] ,
         \decoder/u_input_shifter/w_data_2[2] ,
         \decoder/u_input_shifter/w_data_2[1] ,
         \decoder/u_input_shifter/w_data_2[0] ,
         \decoder/u_input_shifter/w_data_1[15] ,
         \decoder/u_input_shifter/w_data_1[14] ,
         \decoder/u_input_shifter/w_data_1[13] ,
         \decoder/u_input_shifter/w_data_1[12] ,
         \decoder/u_input_shifter/w_data_1[11] ,
         \decoder/u_input_shifter/w_data_1[10] ,
         \decoder/u_input_shifter/w_data_1[9] ,
         \decoder/u_input_shifter/w_data_1[8] ,
         \decoder/u_input_shifter/w_data_1[7] ,
         \decoder/u_input_shifter/w_data_1[6] ,
         \decoder/u_input_shifter/w_data_1[5] ,
         \decoder/u_input_shifter/w_data_1[4] ,
         \decoder/u_input_shifter/w_data_1[3] ,
         \decoder/u_input_shifter/w_data_1[2] ,
         \decoder/u_input_shifter/w_data_1[1] ,
         \decoder/u_input_shifter/w_data_1[0] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_4[2] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_3[2] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_3[3] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_3[4] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_3[5] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_3[6] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_1[2] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_1[3] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_1[4] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_1[5] ,
         \decoder/u_ACS_matrix/w_data_7_to_8_1[6] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_4[3] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_4[4] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_4[5] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_4[6] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_3[0] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_3[1] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_3[2] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_3[3] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_3[4] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_3[5] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_3[6] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_2[0] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_2[1] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_2[4] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_2[5] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_2[6] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_1[0] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_1[1] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_1[2] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_1[3] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_1[4] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_1[5] ,
         \decoder/u_ACS_matrix/w_PM_7_to_8_1[6] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_4[2] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_4[3] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_4[4] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_4[5] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_3[2] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_3[3] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_3[4] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_3[5] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_2[2] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_1[2] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_1[3] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_1[4] ,
         \decoder/u_ACS_matrix/w_data_6_to_7_1[5] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_4[0] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_4[1] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_4[2] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_4[3] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_4[4] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_4[5] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_3[0] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_3[1] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_3[2] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_3[3] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_3[4] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_3[5] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_2[0] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_2[4] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_2[5] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_1[0] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_1[1] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_1[2] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_1[3] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_1[4] ,
         \decoder/u_ACS_matrix/w_PM_6_to_7_1[5] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_4[1] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_4[2] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_4[3] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_4[4] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_3[2] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_3[3] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_3[4] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_2[1] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_2[2] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_2[3] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_2[4] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_1[2] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_1[3] ,
         \decoder/u_ACS_matrix/w_data_5_to_6_1[4] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_4[0] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_4[1] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_4[2] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_4[3] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_4[4] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_3[0] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_3[1] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_3[2] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_3[3] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_3[4] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_2[0] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_2[1] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_2[2] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_2[3] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_2[4] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_1[0] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_1[1] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_1[2] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_1[3] ,
         \decoder/u_ACS_matrix/w_PM_5_to_6_1[4] ,
         \decoder/u_ACS_matrix/w_data_4_to_5_4[2] ,
         \decoder/u_ACS_matrix/w_data_4_to_5_3[2] ,
         \decoder/u_ACS_matrix/w_data_4_to_5_2[2] ,
         \decoder/u_ACS_matrix/w_data_4_to_5_2[3] ,
         \decoder/u_ACS_matrix/w_data_4_to_5_1[2] ,
         \decoder/u_ACS_matrix/w_data_4_to_5_1[3] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_4[0] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_4[2] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_3[0] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_3[1] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_3[2] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_3[3] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_2[0] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_2[1] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_2[2] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_2[3] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_1[0] ,
         \decoder/u_ACS_matrix/w_PM_4_to_5_1[1] ,
         \decoder/u_ACS_matrix/w_data_3_to_4_4[1] ,
         \decoder/u_ACS_matrix/w_data_3_to_4_4[2] ,
         \decoder/u_ACS_matrix/w_data_3_to_4_3[2] ,
         \decoder/u_ACS_matrix/w_data_3_to_4_2[1] ,
         \decoder/u_ACS_matrix/w_data_3_to_4_2[2] ,
         \decoder/u_ACS_matrix/w_data_3_to_4_1[2] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_4[0] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_4[1] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_4[2] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_3[0] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_3[1] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_3[2] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_2[0] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_2[1] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_2[2] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_1[0] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_1[1] ,
         \decoder/u_ACS_matrix/w_PM_3_to_4_1[2] ,
         \decoder/u_ACS_matrix/w_data_2_to_3_2[1] ,
         \decoder/u_ACS_matrix/w_PM_2_to_3_4[0] ,
         \decoder/u_ACS_matrix/w_PM_2_to_3_4[1] ,
         \decoder/u_ACS_matrix/w_PM_2_to_3_3[0] ,
         \decoder/u_ACS_matrix/w_PM_2_to_3_3[1] ,
         \decoder/u_ACS_matrix/w_PM_2_to_3_2[0] ,
         \decoder/u_ACS_matrix/w_PM_2_to_3_2[1] ,
         \decoder/u_ACS_matrix/w_PM_2_to_3_1[0] ,
         \decoder/u_ACS_matrix/w_PM_2_to_3_1[1] ,
         \decoder/u_ACS_matrix/w_PM_1_to_2_4[0] ,
         \decoder/u_ACS_matrix/w_PM_1_to_2_3[0] ,
         \decoder/u_ACS_matrix/w_PM_1_to_2_1[0] , \decoder/u_cmp_sel/N49 ,
         \decoder/u_cmp_sel/N48 , \decoder/u_cmp_sel/N47 ,
         \decoder/u_cmp_sel/N46 , \decoder/u_cmp_sel/N45 ,
         \decoder/u_cmp_sel/N44 , \decoder/u_cmp_sel/N43 ,
         \decoder/u_cmp_sel/N42 ,
         \decoder/u_input_shifter/u_input_fifo/net6035 ,
         \decoder/u_input_shifter/u_input_fifo/net6030 ,
         \decoder/u_input_shifter/u_input_fifo/net6025 ,
         \decoder/u_input_shifter/u_input_fifo/net6020 ,
         \decoder/u_input_shifter/u_input_fifo/net6015 ,
         \decoder/u_input_shifter/u_input_fifo/net6010 ,
         \decoder/u_input_shifter/u_input_fifo/net6005 ,
         \decoder/u_input_shifter/u_input_fifo/net5999 ,
         \decoder/u_input_shifter/u_input_fifo/N28 ,
         \decoder/u_input_shifter/u_input_fifo/N8 ,
         \decoder/u_input_shifter/U_input_split/N51 ,
         \decoder/u_input_shifter/U_input_split/N49 ,
         \decoder/u_input_shifter/U_input_split/N47 ,
         \decoder/u_input_shifter/U_input_split/N45 ,
         \decoder/u_input_shifter/U_input_split/N43 ,
         \decoder/u_input_shifter/U_input_split/N41 ,
         \decoder/u_input_shifter/U_input_split/N39 ,
         \decoder/u_ACS_matrix/u_ACS_col_1/u_ACS_mem_3/u_ACS/ham_dist_2[0] ,
         n311, n313, n315, n317, n318, n320, n322, n324, n326, n328, n330,
         n332, n334, n338, n340, n342, n344, n345, n347, n348, n350, n463,
         n465, n482, n484, n487, n666, n667, n668, n669, n670, n671, n672,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n794,
         n796, n797, n798, n799, n803, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n818, n819, n820, n821, n822, n823, n824, n825,
         n829, n830, n831, n832, n833, n834, n835, n836, n839, n840, n841,
         n842, n843, n844, n845, n846, n850, n851, n852, n853, n854, n855,
         n856, n857, n861, n862, n863, n864, n871, n872, n873, n874, n876,
         n880, n881, n882, n883, n884, n885, n890, n891, n892, n893, n894,
         n895, n900, n901, n902, n903, n909, n910, n911, n912, n917, n918,
         n919, n920, n926, n927, n928, n929, n931, n932, n935, n936, n938,
         n939, n942, n943, n948, n949, n950, n951, n952, n953, n956, n957,
         n958, n959, n960, n961, n963, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1074, n1076, n1080,
         n1082, n1084, n1086, n1088, n1090, n1092, n1094, n1095, n1097, n1098,
         n1100, n1102, n1103, n1108, n1112, n1114, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1144, n1145, n1146, n1147, n1148, n1149, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1323, n1325,
         n1327, n1328, n1330, n1332, n1334, n1336, n1338, n1340, n1342, n1345,
         n1347, n1349, n1351, n1353, n1355, n1357, n1359, n1361, n1363, n1365,
         n1367, n1369, n1371, n1373, n1375, n1377, n1379, n1381, n1383, n1385,
         n1387, n1389, n1391, n1394, n1396, n1400, n1402, n1404, n1406, n1408,
         n1410, n1412, n1414, n1416, n1418, n1420, n1422, n1424, n1426, n1428,
         n1430, n1432, n1433, n1434, n1436, n1438, n1440, n1442, n1444, n1448,
         n1450, n1452, n1454, n1456, n1458, n1460, n1462, n1464, n1466, n1468,
         n1470, n1474, n1476, n1478, n1480, n1482, n1484, n1486, n1488, n1490,
         n1492, n1496, n1498, n1500, n1502, n1505, n1507, n1509, n1511, n1513,
         n1515, n1517, n1519, n1521, n1523, n1525, n1528, n1530, n1532, n1534,
         n1536, n1538, n1540, n1542, n1544, n1546, n1548, n1550, n1552, n1554,
         n1557, n1558, n1559, n1561, n1563, n1565, n1567, n1569, n1571, n1573,
         n1575, n1577, n1579, n1581, n1583, n1585, n1587, n1589, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3032, n3034, n3035, n3036, n3037, n3038, n3039, n3065,
         n3066, n3067, n3068, n3069, n3074, n3076, n3078, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098;
  wire   [15:0] io_data_recv;
  wire   [7:0] io_data_dec;
  tri   clk_PAD;
  tri   rst_PAD;
  tri   [15:0] data_recv_PAD;
  tri   [7:0] data_dec_PAD;

  PDC0204CDG_18 PAD1 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(clk_PAD), .C(io_clk) );
  PDC0204CDG_18 PAD2 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(rst_PAD), .C(io_rst) );
  PDC0204CDG_18 PAD3 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[0]), .C(io_data_recv[0]) );
  PDC0204CDG_18 PAD4 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[1]), .C(io_data_recv[1]) );
  PDC0204CDG_18 PAD5 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[2]), .C(io_data_recv[2]) );
  PDC0204CDG_18 PAD6 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[3]), .C(io_data_recv[3]) );
  PDC0204CDG_18 PAD7 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[4]), .C(io_data_recv[4]) );
  PDC0204CDG_18 PAD8 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[5]), .C(io_data_recv[5]) );
  PDC0204CDG_18 PAD9 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[6]), .C(io_data_recv[6]) );
  PDC0204CDG_18 PAD10 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[7]), .C(io_data_recv[7]) );
  PDC0204CDG_18 PAD11 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[8]), .C(io_data_recv[8]) );
  PDC0204CDG_18 PAD12 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[9]), .C(io_data_recv[9]) );
  PDC0204CDG_18 PAD13 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[10]), .C(io_data_recv[10]) );
  PDC0204CDG_18 PAD14 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[11]), .C(io_data_recv[11]) );
  PDC0204CDG_18 PAD15 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[12]), .C(io_data_recv[12]) );
  PDC0204CDG_18 PAD16 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[13]), .C(io_data_recv[13]) );
  PDC0204CDG_18 PAD17 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[14]), .C(io_data_recv[14]) );
  PDC0204CDG_18 PAD18 ( .I(1'b0), .DS(1'b1), .OEN(1'b1), .PS(1'b0), .PE(1'b0), 
        .IE(1'b1), .PAD(data_recv_PAD[15]), .C(io_data_recv[15]) );
  PDC0204CDG_18 PAD19 ( .I(io_data_dec[0]), .DS(1'b1), .OEN(1'b0), .PS(1'b0), 
        .PE(1'b0), .IE(1'b0), .PAD(data_dec_PAD[0]) );
  PDC0204CDG_18 PAD20 ( .I(io_data_dec[1]), .DS(1'b1), .OEN(1'b0), .PS(1'b0), 
        .PE(1'b0), .IE(1'b0), .PAD(data_dec_PAD[1]) );
  PDC0204CDG_18 PAD21 ( .I(io_data_dec[2]), .DS(1'b1), .OEN(1'b0), .PS(1'b0), 
        .PE(1'b0), .IE(1'b0), .PAD(data_dec_PAD[2]) );
  PDC0204CDG_18 PAD22 ( .I(io_data_dec[3]), .DS(1'b1), .OEN(1'b0), .PS(1'b0), 
        .PE(1'b0), .IE(1'b0), .PAD(data_dec_PAD[3]) );
  PDC0204CDG_18 PAD23 ( .I(io_data_dec[4]), .DS(1'b1), .OEN(1'b0), .PS(1'b0), 
        .PE(1'b0), .IE(1'b0), .PAD(data_dec_PAD[4]) );
  PDC0204CDG_18 PAD24 ( .I(io_data_dec[5]), .DS(1'b1), .OEN(1'b0), .PS(1'b0), 
        .PE(1'b0), .IE(1'b0), .PAD(data_dec_PAD[5]) );
  PDC0204CDG_18 PAD25 ( .I(io_data_dec[6]), .DS(1'b1), .OEN(1'b0), .PS(1'b0), 
        .PE(1'b0), .IE(1'b0), .PAD(data_dec_PAD[6]) );
  PDC0204CDG_18 PAD26 ( .I(io_data_dec[7]), .DS(1'b1), .OEN(1'b0), .PS(1'b0), 
        .PE(1'b0), .IE(1'b0), .PAD(data_dec_PAD[7]) );
  SDFFRHQX2 \decoder/u_input_shifter/U_input_split/out_bit_2_reg[0]  ( .D(
        \decoder/u_input_shifter/U_input_split/N39 ), .SI(1'b0), .SE(1'b0), 
        .CK(io_clk), .RN(n1629), .Q(\decoder/w_enc_bit_2[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_1/u_MEM/PM_out_reg[0]  ( 
        .D(n943), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_PM_2_to_3_1[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_4/u_MEM/PM_out_reg[1]  ( 
        .D(n931), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_PM_2_to_3_4[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_1/u_MEM/PM_out_reg[1]  ( 
        .D(n927), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_1[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_2/u_MEM/PM_out_reg[1]  ( 
        .D(n918), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_2[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_2/u_MEM/PM_out_reg[0]  ( 
        .D(n919), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_2[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_3/u_MEM/PM_out_reg[2]  ( 
        .D(n909), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_3[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_3/u_MEM/PM_out_reg[1]  ( 
        .D(n910), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_3[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_3/u_MEM/PM_out_reg[0]  ( 
        .D(n911), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_3[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_4/u_MEM/PM_out_reg[1]  ( 
        .D(n901), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_4[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_4/u_MEM/PM_out_reg[0]  ( 
        .D(n902), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_4[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_1/u_MEM/PM_out_reg[1]  ( 
        .D(n892), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_1[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_2/u_MEM/PM_out_reg[3]  ( 
        .D(n880), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_2[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_2/u_MEM/PM_out_reg[2]  ( 
        .D(n881), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_2[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_2/u_MEM/PM_out_reg[1]  ( 
        .D(n882), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_2[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_3/u_MEM/PM_out_reg[2]  ( 
        .D(n872), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_3[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_3/u_MEM/PM_out_reg[0]  ( 
        .D(n874), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_3[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_4/u_MEM/PM_out_reg[0]  ( 
        .D(n864), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_4[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_3/u_MEM/PM_out_reg[3]  ( 
        .D(n830), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n3039), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_3[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_3/u_MEM/PM_out_reg[1]  ( 
        .D(n832), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_3[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/PM_out_reg[0]  ( 
        .D(n811), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_1[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/PM_out_reg[2]  ( 
        .D(n786), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_3[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/PM_out_reg[5]  ( 
        .D(n771), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_4[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/PM_out_reg[5]  ( 
        .D(n759), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_2/u_MEM/PM_out_reg[5]  ( 
        .D(n746), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_2[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_2/u_MEM/PM_out_reg[4]  ( 
        .D(n747), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_2[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_2/u_MEM/PM_out_reg[1]  ( 
        .D(n750), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_2[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/PM_out_reg[5]  ( 
        .D(n734), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_1/u_MEM/PM_out_reg[5]  ( 
        .D(n708), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/w_PM_1[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_1/u_MEM/PM_out_reg[0]  ( 
        .D(n713), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/w_PM_1[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_4/u_MEM/PM_out_reg[6]  ( 
        .D(n666), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n3039), .Q(
        \decoder/w_PM_4[6] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_3/u_MEM/PM_out_reg[6]  ( 
        .D(n680), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/w_PM_3[6] ) );
  SDFFSHQX4 R_106 ( .D(n326), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), 
        .Q(n328) );
  SDFFSHQX8 R_2 ( .D(n1591), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n2737) );
  SDFFRHQX8 R_8 ( .D(n1587), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), 
        .Q(n2211) );
  SDFFRQX2 R_10 ( .D(n1822), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), 
        .Q(n1585) );
  SDFFSQXL R_11 ( .D(n1821), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1583) );
  SDFFRQX2 R_14 ( .D(n983), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        n1581) );
  SDFFSQXL R_15 ( .D(n1818), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1579) );
  SDFFSHQX4 R_18 ( .D(n3098), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), 
        .Q(n1575) );
  SDFFSHQX4 R_17 ( .D(n2580), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), 
        .Q(n1577) );
  SDFFSHQX4 R_75 ( .D(n342), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1633), 
        .Q(n344) );
  SDFFSHQX4 R_27 ( .D(n2584), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1629), 
        .Q(n1567) );
  SDFFSHQX4 R_26 ( .D(n2585), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1625), 
        .Q(n1569) );
  SDFFSHQX4 R_33 ( .D(n1557), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1632), 
        .Q(n2175) );
  SDFFRQX2 R_44 ( .D(n2377), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), 
        .Q(n1548) );
  SDFFRHQX8 R_65 ( .D(n1540), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), 
        .Q(n2012) );
  SDFFSHQX2 R_66 ( .D(n2782), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1538) );
  SDFFRHQX4 R_76 ( .D(n1528), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), 
        .Q(n1608) );
  SDFFSHQX4 R_78 ( .D(n2304), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1631), 
        .Q(n1523) );
  SDFFSHQX4 R_77 ( .D(n1328), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1525) );
  SDFFSHQX4 R_83 ( .D(n2791), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), 
        .Q(n1519) );
  SDFFSHQX4 R_96 ( .D(n1174), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1625), 
        .Q(n1505) );
  SDFFSHQX4 R_95 ( .D(n2785), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1632), 
        .Q(n1507) );
  SDFFSHQX8 R_98 ( .D(n334), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1613) );
  SDFFRHQX8 R_105 ( .D(\decoder/u_input_shifter/U_input_split/N43 ), .SI(1'b0), 
        .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(\decoder/w_enc_bit_4[0] ) );
  SDFFRHQX8 R_107 ( .D(n1496), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), 
        .Q(n1897) );
  SDFFSHQX4 R_112 ( .D(n2531), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1625), 
        .Q(n1490) );
  SDFFSHQX4 R_111 ( .D(n2532), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), 
        .Q(n1492) );
  SDFFSHQX4 R_127 ( .D(n2577), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1478) );
  SDFFSHQX4 R_126 ( .D(n3019), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1626), 
        .Q(n1480) );
  SDFFRHQX8 R_159 ( .D(n3037), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), 
        .Q(n1438) );
  SDFFSHQX4 R_186 ( .D(n1927), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1633), 
        .Q(n1402) );
  SDFFSHQX4 R_185 ( .D(n1928), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), 
        .Q(n1404) );
  SDFFRHQX4 R_189 ( .D(\decoder/u_input_shifter/U_input_split/N45 ), .SI(1'b0), 
        .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(\decoder/w_enc_bit_5[0] ) );
  SDFFSHQX4 R_188 ( .D(n330), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), 
        .Q(n332) );
  SDFFSHQX8 R_190 ( .D(n1400), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), 
        .Q(n2011) );
  SDFFSHQX4 R_195 ( .D(n338), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1626), 
        .Q(n1611) );
  SDFFSHQX4 R_197 ( .D(n2708), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), 
        .Q(n1389) );
  SDFFSQXL R_202 ( .D(n2523), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1383) );
  SDFFSHQX4 R_216 ( .D(n1103), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1632), 
        .Q(n1357) );
  SDFFRHQX8 R_220 ( .D(n1355), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), 
        .Q(n2597) );
  SDFFSHQX4 R_222 ( .D(n2704), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1633), 
        .Q(n1351) );
  SDFFSHQX4 R_221 ( .D(n2705), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1631), 
        .Q(n1353) );
  SDFFSQXL R_225 ( .D(n1879), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1347) );
  SDFFSHQX4 R_228 ( .D(n1345), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), 
        .Q(n2210) );
  SDFFSHQX4 R_234 ( .D(n2308), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1632), 
        .Q(n1340) );
  SDFFSHQX4 R_233 ( .D(n2309), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1342) );
  SDFFSHQX4 R_237 ( .D(n2697), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1629), 
        .Q(n1334) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_4/u_MEM/PM_out_reg[2]  ( 
        .D(n820), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_4/u_MEM/PM_out_reg[3]  ( 
        .D(n819), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[3] ) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_2/u_MEM/PM_out_reg[6]  ( 
        .D(n693), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/w_PM_2[6] ) );
  SDFFSHQX2 \decoder/u_input_shifter/U_input_split/out_bit_2_reg[1]  ( .D(n311), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), .Q(n313) );
  SDFFSHQX4 \decoder/u_input_shifter/u_input_fifo/counter_reg[1]  ( .D(n482), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1629), .Q(n484) );
  SDFFRHQX2 R_32 ( .D(n776), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), 
        .Q(\decoder/u_ACS_matrix/w_PM_6_to_7_4[0] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_1/u_MEM/PM_out_reg[0]  ( 
        .D(n854), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_1[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_2/u_MEM/PM_out_reg[1]  ( 
        .D(n842), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_2[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/PM_out_reg[4]  ( 
        .D(n772), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_4[4] ) );
  SDFFSHQX8 \decoder/u_input_shifter/U_input_split/counter_reg[0]  ( .D(n2986), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1633), .Q(n487) );
  SDFFRQX2 R_141 ( .D(1'b1), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), 
        .Q(n1462) );
  SDFFSHQX8 R_5 ( .D(n1589), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), 
        .Q(n2604) );
  SDFFRHQX8 R_25 ( .D(n1571), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), 
        .Q(n2722) );
  SDFFSHQX1 R_58 ( .D(n2788), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1632), 
        .Q(n1542) );
  SDFFSQX2 R_174 ( .D(n2524), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1632), 
        .Q(n1414) );
  SDFFRHQX2 R_227 ( .D(n833), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), 
        .Q(\decoder/u_ACS_matrix/w_PM_5_to_6_3[0] ) );
  SDFFSQXL R_123 ( .D(n1007), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1484) );
  SDFFSQX2 R_135 ( .D(n987), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), 
        .Q(n1470) );
  SDFFSHQX2 R_196 ( .D(n2709), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), 
        .Q(n1391) );
  SDFFSQXL R_212 ( .D(n2517), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1363) );
  SDFFSHQX1 R_84 ( .D(n2790), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1626), 
        .Q(n1517) );
  SDFFSHQX1 R_240 ( .D(n2383), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1625), 
        .Q(n1330) );
  SDFFRHQX4 R_257 ( .D(\decoder/u_input_shifter/U_input_split/N47 ), .SI(1'b0), 
        .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(\decoder/w_enc_bit_6[0] ) );
  SDFFSQXL \decoder/u_input_shifter/U_input_split/out_bit_1_reg[0]  ( .D(n315), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), .Q(n317) );
  SDFFSQX2 R_29 ( .D(n2780), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1563) );
  SDFFSHQX1 R_215 ( .D(n2707), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1633), 
        .Q(n1359) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/PM_out_reg[5]  ( 
        .D(n806), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_1[5] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[13]  ( .D(
        io_data_recv[13]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_4[13] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[12]  ( .D(
        io_data_recv[12]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_4[12] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[9]  ( .D(
        io_data_recv[9]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_4[9] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[8]  ( .D(
        io_data_recv[8]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_4[8] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[7]  ( .D(
        io_data_recv[7]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_4[7] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[4]  ( .D(
        io_data_recv[4]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_4[4] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[1]  ( .D(
        io_data_recv[1]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1625), .Q(
        \decoder/u_input_shifter/w_data_4[1] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[0]  ( .D(
        io_data_recv[0]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_4[0] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[14]  ( .D(
        io_data_recv[14]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_1[14] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[11]  ( .D(
        io_data_recv[11]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_1[11] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[10]  ( .D(
        io_data_recv[10]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_1[10] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[7]  ( .D(
        io_data_recv[7]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_1[7] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[6]  ( .D(
        io_data_recv[6]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_1[6] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[3]  ( .D(
        io_data_recv[3]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_1[3] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[2]  ( .D(
        io_data_recv[2]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_1[2] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[13]  ( .D(
        io_data_recv[13]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_2[13] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[12]  ( .D(
        io_data_recv[12]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_2[12] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[9]  ( .D(
        io_data_recv[9]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_2[9] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[8]  ( .D(
        io_data_recv[8]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_2[8] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[5]  ( .D(
        io_data_recv[5]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_2[5] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[4]  ( .D(
        io_data_recv[4]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_2[4] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[1]  ( .D(
        io_data_recv[1]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_2[1] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[0]  ( .D(
        io_data_recv[0]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_2[0] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[15]  ( .D(
        io_data_recv[15]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_8[15] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[13]  ( .D(
        io_data_recv[13]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_8[13] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[12]  ( .D(
        io_data_recv[12]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1625), .Q(
        \decoder/u_input_shifter/w_data_8[12] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[11]  ( .D(
        io_data_recv[11]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_8[11] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[9]  ( .D(
        io_data_recv[9]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_8[9] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[8]  ( .D(
        io_data_recv[8]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_8[8] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[5]  ( .D(
        io_data_recv[5]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_8[5] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[4]  ( .D(
        io_data_recv[4]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_8[4] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[0]  ( .D(
        io_data_recv[0]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_8[0] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[15]  ( .D(
        io_data_recv[15]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_5[15] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[14]  ( .D(
        io_data_recv[14]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_5[14] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[11]  ( .D(
        io_data_recv[11]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1625), .Q(
        \decoder/u_input_shifter/w_data_5[11] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[10]  ( .D(
        io_data_recv[10]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_5[10] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[7]  ( .D(
        io_data_recv[7]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_5[7] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[6]  ( .D(
        io_data_recv[6]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_5[6] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[5]  ( .D(
        io_data_recv[5]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_5[5] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[3]  ( .D(
        io_data_recv[3]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_5[3] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[2]  ( .D(
        io_data_recv[2]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_5[2] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[1]  ( .D(
        io_data_recv[1]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_5[1] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[15]  ( .D(
        io_data_recv[15]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_6[15] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[13]  ( .D(
        io_data_recv[13]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_6[13] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[12]  ( .D(
        io_data_recv[12]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_6[12] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[9]  ( .D(
        io_data_recv[9]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1625), .Q(
        \decoder/u_input_shifter/w_data_6[9] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[8]  ( .D(
        io_data_recv[8]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_6[8] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[5]  ( .D(
        io_data_recv[5]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_6[5] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[4]  ( .D(
        io_data_recv[4]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_6[4] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[0]  ( .D(
        io_data_recv[0]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_6[0] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[14]  ( .D(
        io_data_recv[14]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_7[14] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[11]  ( .D(
        io_data_recv[11]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_7[11] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[10]  ( .D(
        io_data_recv[10]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_7[10] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[7]  ( .D(
        io_data_recv[7]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1625), .Q(
        \decoder/u_input_shifter/w_data_7[7] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[6]  ( .D(
        io_data_recv[6]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n3039), .Q(
        \decoder/u_input_shifter/w_data_7[6] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[3]  ( .D(
        io_data_recv[3]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n3039), .Q(
        \decoder/u_input_shifter/w_data_7[3] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[2]  ( .D(
        io_data_recv[2]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_7[2] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[1]  ( .D(
        io_data_recv[1]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1625), .Q(
        \decoder/u_input_shifter/w_data_7[1] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[15]  ( .D(
        io_data_recv[15]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_3[15] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[14]  ( .D(
        io_data_recv[14]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_3[14] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[10]  ( .D(
        io_data_recv[10]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_3[10] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[6]  ( .D(
        io_data_recv[6]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_3[6] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[3]  ( .D(
        io_data_recv[3]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_3[3] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[2]  ( .D(
        io_data_recv[2]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_3[2] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[15]  ( .D(
        io_data_recv[15]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_4[15] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[14]  ( .D(
        io_data_recv[14]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_4[14] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[11]  ( .D(
        io_data_recv[11]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_4[11] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[10]  ( .D(
        io_data_recv[10]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_4[10] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[6]  ( .D(
        io_data_recv[6]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_4[6] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[5]  ( .D(
        io_data_recv[5]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_4[5] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[3]  ( .D(
        io_data_recv[3]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_4[3] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_4_reg[2]  ( .D(
        io_data_recv[2]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_4[2] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[15]  ( .D(
        io_data_recv[15]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_1[15] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[13]  ( .D(
        io_data_recv[13]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_1[13] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[12]  ( .D(
        io_data_recv[12]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_1[12] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[9]  ( .D(
        io_data_recv[9]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_1[9] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[8]  ( .D(
        io_data_recv[8]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_1[8] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[5]  ( .D(
        io_data_recv[5]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_1[5] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[4]  ( .D(
        io_data_recv[4]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_1[4] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[1]  ( .D(
        io_data_recv[1]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_1[1] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_1_reg[0]  ( .D(
        io_data_recv[0]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_1[0] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[15]  ( .D(
        io_data_recv[15]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_2[15] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[14]  ( .D(
        io_data_recv[14]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_2[14] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[11]  ( .D(
        io_data_recv[11]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_2[11] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[10]  ( .D(
        io_data_recv[10]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_2[10] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[7]  ( .D(
        io_data_recv[7]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_2[7] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[6]  ( .D(
        io_data_recv[6]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_2[6] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[3]  ( .D(
        io_data_recv[3]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_2[3] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_2_reg[2]  ( .D(
        io_data_recv[2]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_2[2] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[14]  ( .D(
        io_data_recv[14]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_8[14] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[10]  ( .D(
        io_data_recv[10]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_8[10] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[7]  ( .D(
        io_data_recv[7]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_8[7] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[6]  ( .D(
        io_data_recv[6]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_8[6] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[3]  ( .D(
        io_data_recv[3]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_8[3] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[2]  ( .D(
        io_data_recv[2]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_8[2] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_8_reg[1]  ( .D(
        io_data_recv[1]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_8[1] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[13]  ( .D(
        io_data_recv[13]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_5[13] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[12]  ( .D(
        io_data_recv[12]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_5[12] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[9]  ( .D(
        io_data_recv[9]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_5[9] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[8]  ( .D(
        io_data_recv[8]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1625), .Q(
        \decoder/u_input_shifter/w_data_5[8] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[4]  ( .D(
        io_data_recv[4]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_5[4] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_5_reg[0]  ( .D(
        io_data_recv[0]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_5[0] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[14]  ( .D(
        io_data_recv[14]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_6[14] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[11]  ( .D(
        io_data_recv[11]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_6[11] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[10]  ( .D(
        io_data_recv[10]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1626), .Q(
        \decoder/u_input_shifter/w_data_6[10] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[7]  ( .D(
        io_data_recv[7]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_6[7] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[6]  ( .D(
        io_data_recv[6]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1632), .Q(
        \decoder/u_input_shifter/w_data_6[6] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[3]  ( .D(
        io_data_recv[3]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_6[3] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[2]  ( .D(
        io_data_recv[2]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_6[2] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_6_reg[1]  ( .D(
        io_data_recv[1]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .RN(n1625), .Q(
        \decoder/u_input_shifter/w_data_6[1] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[15]  ( .D(
        io_data_recv[15]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_7[15] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[13]  ( .D(
        io_data_recv[13]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_7[13] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[12]  ( .D(
        io_data_recv[12]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_7[12] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[9]  ( .D(
        io_data_recv[9]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_7[9] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[8]  ( .D(
        io_data_recv[8]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_7[8] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[5]  ( .D(
        io_data_recv[5]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1628), .Q(
        \decoder/u_input_shifter/w_data_7[5] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[4]  ( .D(
        io_data_recv[4]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1627), .Q(
        \decoder/u_input_shifter/w_data_7[4] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_7_reg[0]  ( .D(
        io_data_recv[0]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_7[0] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[13]  ( .D(
        io_data_recv[13]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_3[13] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[12]  ( .D(
        io_data_recv[12]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1634), .Q(
        \decoder/u_input_shifter/w_data_3[12] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[11]  ( .D(
        io_data_recv[11]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1635), .Q(
        \decoder/u_input_shifter/w_data_3[11] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[9]  ( .D(
        io_data_recv[9]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1629), .Q(
        \decoder/u_input_shifter/w_data_3[9] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[8]  ( .D(
        io_data_recv[8]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1625), .Q(
        \decoder/u_input_shifter/w_data_3[8] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[7]  ( .D(
        io_data_recv[7]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_3[7] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[5]  ( .D(
        io_data_recv[5]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_3[5] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[4]  ( .D(
        io_data_recv[4]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1630), .Q(
        \decoder/u_input_shifter/w_data_3[4] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[1]  ( .D(
        io_data_recv[1]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1631), .Q(
        \decoder/u_input_shifter/w_data_3[1] ) );
  SDFFRQX2 \decoder/u_input_shifter/u_input_fifo/data_out_3_reg[0]  ( .D(
        io_data_recv[0]), .SI(1'b0), .SE(1'b0), .CK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .RN(n1633), .Q(
        \decoder/u_input_shifter/w_data_3[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_4/u_MEM/PM_out_reg[4]  ( 
        .D(n722), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_4[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/PM_out_reg[1]  ( 
        .D(n810), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_1[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_3/u_MEM/PM_out_reg[2]  ( 
        .D(n831), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_3[2] ) );
  SDFFSQXL \decoder/u_input_shifter/U_input_split/out_bit_1_reg[1]  ( .D(n318), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), .Q(n320) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_1/u_MEM/PM_out_reg[1]  ( 
        .D(n712), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/w_PM_1[1] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_2/u_MEM/PM_out_reg[0]  ( 
        .D(n883), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_2[0] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/data_out_reg[2]  ( 
        .D(n780), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_4[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/PM_out_reg[3]  ( 
        .D(n761), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[3] ) );
  SDFFSHQX4 R_134 ( .D(n1474), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1631), 
        .Q(n1751) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/PM_out_reg[1]  ( 
        .D(n738), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[1] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_3/u_MEM/PM_out_reg[4]  ( 
        .D(n829), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_3[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_1/u_MEM/PM_out_reg[3]  ( 
        .D(n710), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/w_PM_1[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/PM_out_reg[3]  ( 
        .D(n808), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_1[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_1/u_MEM/PM_out_reg[2]  ( 
        .D(n852), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_1[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_2/u_MEM/PM_out_reg[3]  ( 
        .D(n840), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_2[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/PM_out_reg[4]  ( 
        .D(n735), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[4] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/PM_out_reg[4]  ( 
        .D(n784), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_3[4] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/PM_out_reg[5]  ( 
        .D(n783), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_3[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/PM_out_reg[3]  ( 
        .D(n736), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_3/u_MEM/PM_out_reg[3]  ( 
        .D(n871), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_3[3] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_1/u_MEM/PM_out_reg[0]  ( 
        .D(n928), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_1[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/PM_out_reg[3]  ( 
        .D(n785), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_3[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_2/u_MEM/PM_out_reg[2]  ( 
        .D(n841), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_2[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_4/u_MEM/PM_out_reg[5]  ( 
        .D(n721), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_4[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_1/u_MEM/PM_out_reg[0]  ( 
        .D(n893), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_1[0] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_2/u_MEM/data_out_reg[1]  ( 
        .D(n1462), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_data_2_to_3_2[1] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_1/u_MEM/data_out_reg[2]  ( 
        .D(n929), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_data_3_to_4_1[2] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_2/u_MEM/data_out_reg[2]  ( 
        .D(n920), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_data_3_to_4_2[2] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_3/u_MEM/data_out_reg[2]  ( 
        .D(n912), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_data_3_to_4_3[2] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_2/u_MEM/data_out_reg[2]  ( 
        .D(n885), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_data_4_to_5_2[2] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_3/u_MEM/data_out_reg[2]  ( 
        .D(n876), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_data_4_to_5_3[2] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_1/u_MEM/data_out_reg[2]  ( 
        .D(n857), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_1[2] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_2/u_MEM/data_out_reg[2]  ( 
        .D(n846), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_2[2] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_4/u_MEM/data_out_reg[2]  ( 
        .D(n825), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_4[2] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_2/u_MEM/PM_out_reg[6]  ( 
        .D(n745), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_2[6] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_4/u_MEM/data_out_reg[2]  ( 
        .D(n731), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_4[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/PM_out_reg[4]  ( 
        .D(n760), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[4] ) );
  SDFFSQX4 \decoder/u_input_shifter/U_input_split/counter_reg[1]  ( .D(n348), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), .Q(n350) );
  SDFFSQX4 \decoder/u_input_shifter/U_input_split/counter_reg[2]  ( .D(n345), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1631), .Q(n347) );
  SDFFRHQX4 R_133 ( .D(\decoder/u_input_shifter/U_input_split/N41 ), .SI(1'b0), 
        .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(\decoder/w_enc_bit_3[0] ) );
  SDFFSQX2 R_93 ( .D(n2540), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), 
        .Q(n1509) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/PM_out_reg[2]  ( 
        .D(n762), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_3/u_MEM/data_out_reg[3]  ( 
        .D(n691), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/w_data_3[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_3/u_MEM/data_out_reg[4]  ( 
        .D(n690), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/w_data_3[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_3/u_MEM/data_out_reg[5]  ( 
        .D(n689), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/w_data_3[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_3/u_MEM/data_out_reg[6]  ( 
        .D(n688), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/w_data_3[6] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_3/u_MEM/data_out_reg[7]  ( 
        .D(n687), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/w_data_3[7] ) );
  SDFFSHQX2 R_165 ( .D(n1119), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), 
        .Q(n1426) );
  SDFFSHQX2 R_164 ( .D(n2543), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), 
        .Q(n1428) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/data_out_reg[3]  ( 
        .D(n768), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_1[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/data_out_reg[6]  ( 
        .D(n765), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_1[6] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/data_out_reg[5]  ( 
        .D(n766), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_1[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/data_out_reg[4]  ( 
        .D(n767), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_1[4] ) );
  SDFFSQX2 R_192 ( .D(n2526), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1633), 
        .Q(n1394) );
  SDFFSHQX8 R_158 ( .D(n2797), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1629), 
        .Q(n1440) );
  SDFFRHQX2 \decoder/u_cmp_sel/data_out_reg[6]  ( .D(\decoder/u_cmp_sel/N48 ), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(io_data_dec[6]) );
  SDFFSHQX4 R_191 ( .D(n1139), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), 
        .Q(n1396) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/data_out_reg[5]  ( 
        .D(n741), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_3[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/data_out_reg[3]  ( 
        .D(n743), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_3[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/data_out_reg[6]  ( 
        .D(n740), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_3[6] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/data_out_reg[4]  ( 
        .D(n742), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_3[4] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_2/u_MEM/data_out_reg[2]  ( 
        .D(n803), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_2[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_2/u_MEM/data_out_reg[4]  ( 
        .D(n844), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n3039), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_2[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_2/u_MEM/data_out_reg[3]  ( 
        .D(n845), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_2[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/data_out_reg[3]  ( 
        .D(n814), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n3039), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_1[3] ) );
  SDFFRHQX4 \decoder/u_cmp_sel/data_out_reg[0]  ( .D(\decoder/u_cmp_sel/N42 ), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(io_data_dec[0]) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_3/u_MEM/data_out_reg[2]  ( 
        .D(n692), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/w_data_3[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/data_out_reg[5]  ( 
        .D(n812), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_1[5] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/data_out_reg[2]  ( 
        .D(n792), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_3[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_1/u_MEM/data_out_reg[3]  ( 
        .D(n894), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_data_4_to_5_1[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_3/u_MEM/data_out_reg[4]  ( 
        .D(n834), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_3[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_3/u_MEM/data_out_reg[3]  ( 
        .D(n835), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_3[3] ) );
  SDFFSHQX4 R_79 ( .D(n2964), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), 
        .Q(n1521) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/PM_out_reg[1]  ( 
        .D(n775), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_4[1] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/PM_out_reg[1]  ( 
        .D(n763), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/data_out_reg[4]  ( 
        .D(n813), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_1[4] ) );
  SDFFRHQX2 \decoder/u_cmp_sel/data_out_reg[7]  ( .D(\decoder/u_cmp_sel/N49 ), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(io_data_dec[7]) );
  SDFFRHQX2 \decoder/u_cmp_sel/data_out_reg[4]  ( .D(\decoder/u_cmp_sel/N46 ), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(io_data_dec[4]) );
  SDFFRHQX2 \decoder/u_cmp_sel/data_out_reg[5]  ( .D(\decoder/u_cmp_sel/N47 ), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(io_data_dec[5]) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_4/u_MEM/data_out_reg[4]  ( 
        .D(n823), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_4[4] ) );
  SDFFSHQX4 R_253 ( .D(n338), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), 
        .Q(n340) );
  SDFFSHQX4 R_256 ( .D(n1108), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1255) );
  SDFFRHQX8 R_258 ( .D(\decoder/u_input_shifter/U_input_split/N47 ), .SI(1'b0), 
        .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(n1248) );
  SDFFSHQX8 R_283 ( .D(n1624), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1631), 
        .Q(n1102) );
  SDFFSHQX8 R_284 ( .D(n3092), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1631), 
        .Q(n1100) );
  SDFFSQXL R_290 ( .D(n2985), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n3039), 
        .Q(n1090) );
  SDFFRQX2 R_291 ( .D(n1820), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), 
        .Q(n1088) );
  SDFFSHQX4 R_132 ( .D(n322), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), 
        .Q(n324) );
  SDFFSQX2 \decoder/u_input_shifter/u_input_fifo/counter_reg[2]  ( .D(n463), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), .Q(n465) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_1/u_MEM/PM_out_reg[6]  ( 
        .D(n707), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/w_PM_1[6] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/data_out_reg[5]  ( 
        .D(n789), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_3[5] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/data_out_reg[4]  ( 
        .D(n790), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_3[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/data_out_reg[3]  ( 
        .D(n791), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_3[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_1/u_MEM/PM_out_reg[4]  ( 
        .D(n850), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_1[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_2/u_MEM/data_out_reg[2]  ( 
        .D(n705), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/w_data_2[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_1/u_MEM/data_out_reg[4]  ( 
        .D(n855), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_1[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_1/u_MEM/data_out_reg[3]  ( 
        .D(n856), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_1[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_2/u_MEM/data_out_reg[3]  ( 
        .D(n884), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_data_4_to_5_2[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_4/u_MEM/data_out_reg[3]  ( 
        .D(n824), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_4[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_2/u_MEM/PM_out_reg[2]  ( 
        .D(n917), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_2[2] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_1/u_MEM/PM_out_reg[3]  ( 
        .D(n851), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_1[3] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/PM_out_reg[3]  ( 
        .D(n773), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_4[3] ) );
  SDFFSHQX4 R_292 ( .D(n2787), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), 
        .Q(n1086) );
  SDFFSHQX4 R_293 ( .D(n3022), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1084) );
  SDFFSHQX2 R_295 ( .D(n1013), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), 
        .Q(n1080) );
  SDFFSHQX8 R_294 ( .D(n2400), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), 
        .Q(n1082) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_2/u_MEM/PM_out_reg[0]  ( 
        .D(n751), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_2[0] ) );
  SDFFRHQX8 R_252 ( .D(\decoder/u_input_shifter/U_input_split/N49 ), .SI(1'b0), 
        .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(\decoder/w_enc_bit_7[0] ) );
  SDFFSHQX2 R_173 ( .D(n2525), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), 
        .Q(n1416) );
  SDFFRHQX2 \decoder/u_cmp_sel/data_out_reg[2]  ( .D(\decoder/u_cmp_sel/N44 ), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(io_data_dec[2]) );
  SDFFSHQX8 R_19 ( .D(n1127), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1626), 
        .Q(n1573) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_2/u_MEM/PM_out_reg[0]  ( 
        .D(n799), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_2[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_1/u_MEM/PM_out_reg[1]  ( 
        .D(n853), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_1[1] ) );
  SDFFSHQX4 R_35 ( .D(n1017), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1625), 
        .Q(n1552) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_2/u_MEM/PM_out_reg[4]  ( 
        .D(n1114), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n3039), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_2[4] ) );
  SDFFSHQX4 R_104 ( .D(n2964), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1629), 
        .Q(n1498) );
  SDFFSHQX2 R_246 ( .D(n2964), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1632), 
        .Q(n1327) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_4/u_MEM/PM_out_reg[1]  ( 
        .D(n821), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_3/u_MEM/PM_out_reg[1]  ( 
        .D(n873), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_3[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_2/u_MEM/PM_out_reg[5]  ( 
        .D(n694), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/w_PM_2[5] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_1/u_MEM/data_out_reg[2]  ( 
        .D(n895), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(
        \decoder/u_ACS_matrix/w_data_4_to_5_1[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/data_out_reg[3]  ( 
        .D(n779), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_4[3] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/data_out_reg[4]  ( 
        .D(n778), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_4[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/data_out_reg[5]  ( 
        .D(n777), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_4[5] ) );
  SDFFSHQX4 R_34 ( .D(n3029), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1626), 
        .Q(n1554) );
  CLKINVX3 U1102 ( .A(n2351), .Y(n2403) );
  DLY1X1 U1103 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_1[1] ), .Y(n956) );
  INVX6 U1106 ( .A(n1158), .Y(n961) );
  NAND2X8 U1107 ( .A(\decoder/w_enc_bit_7[0] ), .B(n340), .Y(n2172) );
  NOR2X4 U1110 ( .A(n958), .B(n2385), .Y(n2185) );
  AOI21X6 U1111 ( .A0(n2203), .A1(n2189), .B0(n2383), .Y(n1262) );
  NOR2X8 U1112 ( .A(n1152), .B(n2176), .Y(n2203) );
  NAND2BX4 U1113 ( .AN(n2411), .B(n2412), .Y(n2344) );
  OR2X4 U1115 ( .A(n2444), .B(n2711), .Y(n1605) );
  INVX10 U1116 ( .A(n2484), .Y(n1019) );
  INVX4 U1119 ( .A(n2405), .Y(n1195) );
  XNOR2X4 U1120 ( .A(n2349), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_2[5] ), .Y(
        n2351) );
  OAI21BX4 U1123 ( .A0(n2363), .A1(\decoder/u_ACS_matrix/w_PM_6_to_7_1[4] ), 
        .B0N(n960), .Y(n2406) );
  XNOR2X4 U1124 ( .A(n960), .B(n959), .Y(n2404) );
  CLKINVX16 U1125 ( .A(n2593), .Y(n959) );
  NAND2X8 U1127 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_4[2] ), .B(
        \decoder/u_ACS_matrix/w_PM_6_to_7_4[1] ), .Y(n2167) );
  AOI31X2 U1129 ( .A0(n957), .A1(n2356), .A2(n2357), .B0(n2407), .Y(n2359) );
  OAI21X8 U1130 ( .A0(n2557), .A1(\decoder/u_ACS_matrix/w_PM_6_to_7_3[0] ), 
        .B0(\decoder/u_ACS_matrix/w_PM_6_to_7_3[1] ), .Y(n2170) );
  OAI211X4 U1131 ( .A0(n2605), .A1(n998), .B0(n2344), .C0(n2614), .Y(n2360) );
  CLKNAND2X12 U1133 ( .A(n961), .B(n1287), .Y(n2955) );
  NAND2X4 U1136 ( .A(n1892), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_2[1] ), .Y(
        n1909) );
  OAI21BX4 U1138 ( .A0(n1750), .A1(n1749), .B0N(n1748), .Y(n1834) );
  OR2X4 U1140 ( .A(n2103), .B(n2100), .Y(n963) );
  NOR2BX8 U1141 ( .AN(n1751), .B(n1708), .Y(n1707) );
  INVX6 U1142 ( .A(n1707), .Y(n1713) );
  INVX2 U1144 ( .A(n833), .Y(n1345) );
  XOR2X2 U1145 ( .A(\decoder/u_ACS_matrix/w_PM_4_to_5_3[3] ), .B(n966), .Y(
        n1977) );
  NAND2BX4 U1147 ( .AN(n1785), .B(n1784), .Y(n1759) );
  OAI21X2 U1148 ( .A0(n1756), .A1(\decoder/u_ACS_matrix/w_PM_2_to_3_2[1] ), 
        .B0(n1754), .Y(n1785) );
  OAI2B11X4 U1149 ( .A1N(n1754), .A0(n1763), .B0(n1762), .C0(n1039), .Y(n1782)
         );
  AOI21X4 U1150 ( .A0(n2050), .A1(n2042), .B0(n1931), .Y(n1937) );
  NAND2X8 U1151 ( .A(n1932), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_4[0] ), .Y(
        n2050) );
  OAI21X2 U1155 ( .A0(\decoder/u_ACS_matrix/w_PM_1_to_2_4[0] ), .A1(n1667), 
        .B0(n1697), .Y(n1701) );
  NAND2X4 U1156 ( .A(n1667), .B(\decoder/u_ACS_matrix/w_PM_1_to_2_4[0] ), .Y(
        n1697) );
  NOR2X4 U1157 ( .A(n1663), .B(n1662), .Y(n1681) );
  NOR2XL U1158 ( .A(n1692), .B(n1694), .Y(n1662) );
  INVXL U1159 ( .A(n2147), .Y(n2149) );
  AND2X6 U1160 ( .A(n2046), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_3[1] ), .Y(
        n2048) );
  NOR2XL U1165 ( .A(n1133), .B(n1938), .Y(n967) );
  AND3X4 U1167 ( .A(n2046), .B(n968), .C(
        \decoder/u_ACS_matrix/w_PM_4_to_5_3[1] ), .Y(n2056) );
  CLKINVX3 U1169 ( .A(n2059), .Y(n969) );
  OAI2BB1X2 U1171 ( .A0N(n1894), .A1N(n1895), .B0(n1896), .Y(n970) );
  BUFX2 U1172 ( .A(n1797), .Y(n971) );
  OAI21X4 U1173 ( .A0(n1770), .A1(\decoder/u_ACS_matrix/w_PM_2_to_3_3[1] ), 
        .B0(n1771), .Y(n1795) );
  NAND2X4 U1177 ( .A(n1920), .B(n976), .Y(n1896) );
  NAND2X4 U1178 ( .A(n2991), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_1[0] ), .Y(
        n1895) );
  OAI21X4 U1179 ( .A0(n1709), .A1(\decoder/u_ACS_matrix/w_PM_2_to_3_2[1] ), 
        .B0(n1715), .Y(n1727) );
  NAND2X4 U1180 ( .A(n1709), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_2[1] ), .Y(
        n1715) );
  NAND2X4 U1181 ( .A(n1753), .B(n1751), .Y(n1709) );
  OR2X4 U1183 ( .A(n1795), .B(n1794), .Y(n1225) );
  OAI21X2 U1184 ( .A0(n2056), .A1(\decoder/u_ACS_matrix/w_PM_4_to_5_3[3] ), 
        .B0(n2099), .Y(n2095) );
  OAI21X2 U1185 ( .A0(n2099), .A1(n2097), .B0(n2064), .Y(n2070) );
  NAND2X8 U1186 ( .A(n2012), .B(n2011), .Y(n1932) );
  OAI2BB1X4 U1187 ( .A0N(n2837), .A1N(n2836), .B0(n2846), .Y(n2838) );
  OAI211X2 U1188 ( .A0(\decoder/w_PM_2[6] ), .A1(n2895), .B0(n2848), .C0(n2847), .Y(n2859) );
  INVX4 U1190 ( .A(n2095), .Y(n2059) );
  NAND2BX8 U1192 ( .AN(n1998), .B(n1183), .Y(n2007) );
  NAND3BX4 U1193 ( .AN(n972), .B(n2055), .C(n2054), .Y(n2060) );
  NOR2X2 U1194 ( .A(n2092), .B(n2090), .Y(n972) );
  OAI2BB1X2 U1195 ( .A0N(n1992), .A1N(n1274), .B0(n2995), .Y(n2144) );
  NAND2BX4 U1197 ( .AN(n2724), .B(n3081), .Y(n973) );
  NAND2BX8 U1198 ( .AN(n2722), .B(n726), .Y(n2732) );
  OAI21X2 U1199 ( .A0(n2044), .A1(n2066), .B0(n863), .Y(n2049) );
  INVXL U1200 ( .A(n979), .Y(n980) );
  INVXL U1202 ( .A(n1279), .Y(n974) );
  NAND2X4 U1207 ( .A(n1839), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_2[3] ), .Y(
        n1861) );
  XNOR2X2 U1208 ( .A(n1998), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_3[2] ), .Y(
        n2143) );
  NAND2BX4 U1209 ( .AN(n2066), .B(n2043), .Y(n1939) );
  INVX4 U1212 ( .A(n2991), .Y(n976) );
  NAND2BX4 U1214 ( .AN(n977), .B(n2654), .Y(n2574) );
  XNOR2X2 U1215 ( .A(n1598), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[5] ), .Y(
        n977) );
  NOR2X2 U1217 ( .A(n2919), .B(n1780), .Y(n903) );
  OAI21X6 U1218 ( .A0(n1691), .A1(n1722), .B0(n1723), .Y(n2919) );
  AOI21X4 U1219 ( .A0(n1871), .A1(n1870), .B0(n1875), .Y(n1922) );
  NAND2X4 U1220 ( .A(n1866), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_4[1] ), .Y(
        n1870) );
  NOR2X8 U1221 ( .A(n1870), .B(n1871), .Y(n1875) );
  AOI2B1X2 U1222 ( .A1N(\decoder/u_ACS_matrix/w_PM_4_to_5_3[2] ), .A0(n1938), 
        .B0(n1935), .Y(n1980) );
  BUFX10 U1223 ( .A(n1092), .Y(n978) );
  OAI2BB1X4 U1225 ( .A0N(n1987), .A1N(n1986), .B0(n1989), .Y(n2160) );
  NAND2BX4 U1226 ( .AN(n1986), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_4[4] ), 
        .Y(n1989) );
  INVXL U1227 ( .A(n2092), .Y(n979) );
  DLY1X1 U1228 ( .A(n980), .Y(n1153) );
  BUFX2 U1229 ( .A(n863), .Y(n981) );
  NOR2X4 U1230 ( .A(n2700), .B(n2699), .Y(n2692) );
  XNOR2X2 U1233 ( .A(n2679), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_4[5] ), .Y(
        n2699) );
  AOI21X2 U1236 ( .A0(n1910), .A1(n1914), .B0(n1190), .Y(n1911) );
  INVX2 U1237 ( .A(n1817), .Y(n983) );
  CLKINVX3 U1239 ( .A(n1869), .Y(n1880) );
  NAND3X4 U1240 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_3[2] ), .B(n1867), .C(
        \decoder/u_ACS_matrix/w_PM_3_to_4_3[1] ), .Y(n1869) );
  NAND2X4 U1241 ( .A(n2096), .B(n2059), .Y(n2064) );
  OAI21X2 U1242 ( .A0(n1934), .A1(n861), .B0(n1933), .Y(n1979) );
  OAI21X4 U1243 ( .A0(n1926), .A1(n1928), .B0(n1873), .Y(n1881) );
  NAND2X4 U1244 ( .A(n1925), .B(n1872), .Y(n1873) );
  OAI211X2 U1245 ( .A0(n1864), .A1(n1874), .B0(n1741), .C0(n1740), .Y(n1745)
         );
  INVX4 U1246 ( .A(n2993), .Y(n1845) );
  NAND2XL U1249 ( .A(n2027), .B(n2082), .Y(n2020) );
  BUFX2 U1254 ( .A(n2224), .Y(n984) );
  NAND2X4 U1256 ( .A(n2644), .B(n2618), .Y(n2609) );
  NAND2X4 U1257 ( .A(n2591), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_1[4] ), .Y(
        n1607) );
  OAI21X2 U1259 ( .A0(n1999), .A1(\decoder/u_ACS_matrix/w_PM_5_to_6_3[1] ), 
        .B0(n1998), .Y(n2142) );
  NOR2XL U1261 ( .A(n2141), .B(n2142), .Y(n2000) );
  INVXL U1262 ( .A(n2033), .Y(n2084) );
  MXI2X1 U1266 ( .A(n2649), .B(n3094), .S0(n1623), .Y(n738) );
  XNOR2X4 U1269 ( .A(n1993), .B(n1990), .Y(n2145) );
  INVX4 U1271 ( .A(n2613), .Y(n985) );
  INVXL U1272 ( .A(n2613), .Y(n2657) );
  NOR2X4 U1273 ( .A(n1851), .B(n2018), .Y(n1839) );
  AOI21X4 U1274 ( .A0(n1957), .A1(n1181), .B0(n1840), .Y(n1858) );
  NOR2X2 U1276 ( .A(n1998), .B(n2218), .Y(n1991) );
  OAI2BB1X2 U1277 ( .A0N(n2003), .A1N(n2002), .B0(n2001), .Y(n2005) );
  NAND2BX4 U1278 ( .AN(n2535), .B(n987), .Y(n2502) );
  NAND3BX2 U1279 ( .AN(n2213), .B(n1313), .C(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[4] ), .Y(n2215) );
  NOR2BX2 U1280 ( .AN(n1313), .B(n2213), .Y(n2242) );
  NAND3X2 U1281 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_4[2] ), .B(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[1] ), .C(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[3] ), .Y(n2213) );
  INVX6 U1282 ( .A(n2483), .Y(n2481) );
  OAI21X2 U1285 ( .A0(n1839), .A1(\decoder/u_ACS_matrix/w_PM_4_to_5_2[3] ), 
        .B0(n1861), .Y(n1961) );
  NAND2X4 U1288 ( .A(n2601), .B(n797), .Y(n2606) );
  NAND3X4 U1289 ( .A(n2235), .B(n2236), .C(n2234), .Y(n2244) );
  INVX2 U1290 ( .A(n2527), .Y(n1123) );
  OAI21X2 U1291 ( .A0(n1599), .A1(\decoder/u_ACS_matrix/w_PM_7_to_8_2[1] ), 
        .B0(n2483), .Y(n2527) );
  NAND3X4 U1292 ( .A(n2495), .B(n2494), .C(n2493), .Y(n2501) );
  NOR2BX4 U1293 ( .AN(n2627), .B(n2655), .Y(n2625) );
  INVX8 U1294 ( .A(n1956), .Y(n1958) );
  INVX4 U1295 ( .A(n863), .Y(n1931) );
  NAND2X4 U1298 ( .A(n1756), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_2[1] ), .Y(
        n1754) );
  OAI211X4 U1299 ( .A0(n1761), .A1(n1760), .B0(n1759), .C0(n1758), .Y(n1762)
         );
  NAND2X2 U1301 ( .A(n2636), .B(n2655), .Y(n1011) );
  NAND2X4 U1302 ( .A(n985), .B(n2592), .Y(n2636) );
  NAND2X4 U1303 ( .A(n2596), .B(n1607), .Y(n2641) );
  NAND2BX4 U1304 ( .AN(n2642), .B(n2641), .Y(n2626) );
  NAND2X2 U1308 ( .A(n2603), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_1[2] ), .Y(
        n2608) );
  NAND2X4 U1309 ( .A(n1592), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_3[4] ), .Y(
        n2165) );
  CLKINVX3 U1310 ( .A(n2007), .Y(n1592) );
  CLKINVX3 U1311 ( .A(n1988), .Y(n2164) );
  OAI21X1 U1313 ( .A0(n1124), .A1(n1144), .B0(n1307), .Y(n987) );
  NAND2X4 U1316 ( .A(n2221), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_4[2] ), .Y(
        n2241) );
  NAND3X4 U1317 ( .A(n2768), .B(n2767), .C(n2775), .Y(n2778) );
  NAND4X8 U1322 ( .A(n989), .B(n2832), .C(n2831), .D(n2830), .Y(n2916) );
  AND4X2 U1323 ( .A(n2802), .B(n2801), .C(n2856), .D(n2800), .Y(n989) );
  NAND2X4 U1325 ( .A(n2164), .B(n2165), .Y(n2161) );
  INVX4 U1326 ( .A(n2573), .Y(n2654) );
  MXI2X2 U1330 ( .A(n1353), .B(n1351), .S0(n1102), .Y(n696) );
  OAI21X2 U1332 ( .A0(n2081), .A1(n2078), .B0(n2020), .Y(n2035) );
  OAI21X2 U1333 ( .A0(n2633), .A1(n2623), .B0(n2631), .Y(n2624) );
  OR2X4 U1334 ( .A(n2606), .B(n1022), .Y(n2595) );
  NAND3BX4 U1336 ( .AN(n2819), .B(n2818), .C(n2820), .Y(n2862) );
  NAND3BX4 U1337 ( .AN(n672), .B(n2817), .C(n686), .Y(n2818) );
  INVX4 U1340 ( .A(n684), .Y(n2824) );
  MXI2X4 U1341 ( .A(n1511), .B(n1509), .S0(n1100), .Y(n684) );
  OAI211X2 U1342 ( .A0(n1966), .A1(n1964), .B0(n1848), .C0(n1847), .Y(n1853)
         );
  AOI2BB2X2 U1343 ( .B0(n2982), .B1(n700), .A0N(n992), .A1N(n993), .Y(n2918)
         );
  INVX12 U1344 ( .A(n1118), .Y(n1145) );
  NAND2X2 U1345 ( .A(n2630), .B(n2629), .Y(n2632) );
  NAND2X8 U1346 ( .A(n2075), .B(n2098), .Y(n2953) );
  OAI21X2 U1347 ( .A0(n2720), .A1(n726), .B0(n2732), .Y(n2786) );
  INVXL U1351 ( .A(n2306), .Y(n2233) );
  NAND2X4 U1352 ( .A(n2420), .B(n2542), .Y(n2421) );
  NAND2BX8 U1354 ( .AN(n2170), .B(n2169), .Y(n994) );
  NAND2X4 U1356 ( .A(n2558), .B(n2579), .Y(n2560) );
  NOR2X4 U1358 ( .A(n2534), .B(n2455), .Y(n2447) );
  OAI21X2 U1359 ( .A0(n2989), .A1(n2481), .B0(n2480), .Y(n2541) );
  NAND2X4 U1360 ( .A(n2989), .B(n2481), .Y(n2480) );
  NAND3X4 U1361 ( .A(n1270), .B(n1269), .C(n2560), .Y(n1130) );
  NAND3X2 U1362 ( .A(n995), .B(n2625), .C(n2624), .Y(n2639) );
  INVXL U1364 ( .A(n2530), .Y(n996) );
  INVX2 U1365 ( .A(n996), .Y(n997) );
  AOI22X2 U1366 ( .A0(n2982), .A1(\decoder/w_data_2[2] ), .B0(n1145), .B1(
        n1071), .Y(n2979) );
  INVX4 U1368 ( .A(n696), .Y(n2869) );
  NOR2X2 U1372 ( .A(n2745), .B(n2779), .Y(n1027) );
  AND4X4 U1373 ( .A(n2725), .B(n1203), .C(n2726), .D(n1201), .Y(n2745) );
  BUFX2 U1374 ( .A(n1235), .Y(n998) );
  NAND2X4 U1376 ( .A(n2200), .B(n1130), .Y(n2192) );
  NAND2X4 U1378 ( .A(n2264), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[1] ), .Y(
        n2271) );
  AOI21X2 U1379 ( .A0(n2273), .A1(n2315), .B0(n2317), .Y(n2279) );
  CLKINVX3 U1380 ( .A(n2181), .Y(n1295) );
  AO21X4 U1381 ( .A0(n2812), .A1(n2811), .B0(n2810), .Y(n2813) );
  AOI21X4 U1382 ( .A0(n2455), .A1(n2456), .B0(n1007), .Y(n2458) );
  OAI21X2 U1383 ( .A0(n3067), .A1(\decoder/u_ACS_matrix/w_PM_7_to_8_2[0] ), 
        .B0(n2471), .Y(n2525) );
  AOI2B1X4 U1384 ( .A1N(n2443), .A0(n2440), .B0(n2439), .Y(n2441) );
  OAI21X2 U1388 ( .A0(n796), .A1(n2345), .B0(n2346), .Y(n2407) );
  NAND3X6 U1389 ( .A(n1019), .B(n1289), .C(n1288), .Y(n2416) );
  NAND2BX4 U1390 ( .AN(\decoder/u_ACS_matrix/w_PM_7_to_8_1[0] ), .B(n2432), 
        .Y(n1289) );
  NOR2BX4 U1391 ( .AN(n2444), .B(n2456), .Y(n2454) );
  INVX4 U1392 ( .A(n698), .Y(n1121) );
  MXI2X2 U1394 ( .A(n1391), .B(n1389), .S0(n1102), .Y(n698) );
  NAND2X2 U1395 ( .A(n1195), .B(n2406), .Y(n999) );
  OAI21X8 U1396 ( .A0(n2340), .A1(n2329), .B0(n1235), .Y(n1010) );
  OAI31X4 U1397 ( .A0(n2844), .A1(n2843), .A2(n2842), .B0(n2841), .Y(n2848) );
  BUFX2 U1398 ( .A(n2546), .Y(n1000) );
  XNOR2X4 U1399 ( .A(n1001), .B(n748), .Y(n2420) );
  XNOR2X4 U1400 ( .A(n1001), .B(n2437), .Y(n2539) );
  NAND2X2 U1401 ( .A(n2417), .B(n1257), .Y(n1001) );
  MXI2X2 U1402 ( .A(n1359), .B(n1357), .S0(n1102), .Y(n697) );
  NAND2X2 U1403 ( .A(n1002), .B(\decoder/w_PM_1[5] ), .Y(n2894) );
  MXI2X6 U1405 ( .A(n1507), .B(n1505), .S0(n1433), .Y(n667) );
  NAND2X8 U1406 ( .A(n1438), .B(n1440), .Y(n1433) );
  INVX4 U1407 ( .A(n2711), .Y(n2455) );
  NOR2X4 U1408 ( .A(n2443), .B(n2442), .Y(n2456) );
  NAND2X4 U1409 ( .A(n2862), .B(n2861), .Y(n2877) );
  NOR2BX4 U1411 ( .AN(n2410), .B(n2409), .Y(n2361) );
  AOI2BB2X2 U1413 ( .B0(n2982), .B1(n704), .A0N(n992), .A1N(n1003), .Y(n2973)
         );
  NAND2X4 U1415 ( .A(\decoder/w_enc_bit_5[0] ), .B(n332), .Y(n2042) );
  NOR2X2 U1417 ( .A(n2070), .B(n2069), .Y(n2071) );
  NAND2X4 U1418 ( .A(n2056), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_3[3] ), .Y(
        n2099) );
  BUFX12 U1419 ( .A(n2597), .Y(n1235) );
  OR2X4 U1420 ( .A(n2521), .B(n2520), .Y(n1004) );
  INVXL U1422 ( .A(n2498), .Y(n1005) );
  INVX2 U1424 ( .A(n2541), .Y(n2498) );
  NAND2X6 U1426 ( .A(n2784), .B(n2766), .Y(n2775) );
  NAND2X4 U1427 ( .A(n2255), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[0] ), .Y(
        n2251) );
  INVXL U1428 ( .A(n2435), .Y(n1006) );
  INVX4 U1429 ( .A(n2542), .Y(n2435) );
  BUFX4 U1430 ( .A(n2712), .Y(n1007) );
  INVXL U1431 ( .A(n2317), .Y(n1008) );
  INVX2 U1432 ( .A(n1008), .Y(n1009) );
  NAND2X4 U1433 ( .A(n2423), .B(n1144), .Y(n2422) );
  INVX4 U1434 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_2[0] ), .Y(n2329) );
  AOI21X4 U1435 ( .A0(n2368), .A1(n2408), .B0(n2367), .Y(n2369) );
  NAND2X4 U1436 ( .A(n2637), .B(n1012), .Y(n2638) );
  INVX2 U1437 ( .A(n1011), .Y(n1012) );
  OR2X4 U1438 ( .A(n1607), .B(n2593), .Y(n2655) );
  NAND2BX4 U1439 ( .AN(n2603), .B(n2600), .Y(n2648) );
  BUFX2 U1441 ( .A(n2710), .Y(n1013) );
  AOI21X2 U1442 ( .A0(n1155), .A1(n2587), .B0(n2586), .Y(n1014) );
  INVX4 U1443 ( .A(n2620), .Y(n2644) );
  INVX2 U1445 ( .A(n2780), .Y(n1016) );
  INVXL U1447 ( .A(n2176), .Y(n1017) );
  NOR2XL U1448 ( .A(n2318), .B(n2274), .Y(n1018) );
  INVX4 U1449 ( .A(n2459), .Y(n2534) );
  XNOR2X4 U1450 ( .A(n2461), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_2[5] ), .Y(
        n2459) );
  NOR2BX4 U1452 ( .AN(n1155), .B(n1189), .Y(n1247) );
  XNOR2X4 U1453 ( .A(n2595), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_2[5] ), .Y(
        n2613) );
  INVX4 U1454 ( .A(n2432), .Y(n2488) );
  NAND3X4 U1455 ( .A(n1206), .B(n2740), .C(n2739), .Y(n2747) );
  NAND2X2 U1456 ( .A(n2741), .B(n2789), .Y(n1206) );
  XNOR2X4 U1457 ( .A(n2174), .B(n1316), .Y(n1251) );
  INVX2 U1459 ( .A(n3010), .Y(n1020) );
  CLKINVX3 U1460 ( .A(n2903), .Y(n2905) );
  OAI2BB1X2 U1463 ( .A0N(n1128), .A1N(n2586), .B0(n2334), .Y(n1024) );
  AOI21X2 U1464 ( .A0(n2622), .A1(n2642), .B0(n2621), .Y(n2631) );
  INVXL U1465 ( .A(n1251), .Y(n2387) );
  NAND2BX4 U1466 ( .AN(n2712), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_2[5] ), 
        .Y(n2439) );
  CLKINVX3 U1472 ( .A(n2406), .Y(n2358) );
  NOR2X4 U1473 ( .A(n2451), .B(n2450), .Y(n2449) );
  NAND2BX2 U1475 ( .AN(n2546), .B(n2545), .Y(n2556) );
  OAI21X4 U1477 ( .A0(n1014), .A1(n797), .B0(n2606), .Y(n2646) );
  OAI2BB1X4 U1478 ( .A0N(n2252), .A1N(n2253), .B0(n2271), .Y(n2321) );
  NAND2X4 U1480 ( .A(n1220), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_2[1] ), .Y(
        n2483) );
  NOR2X4 U1482 ( .A(n2190), .B(n2547), .Y(n2194) );
  XNOR2X2 U1483 ( .A(n2194), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[5] ), .Y(
        n2379) );
  MXI2X2 U1484 ( .A(n1086), .B(n1084), .S0(n1433), .Y(n672) );
  OAI21X1 U1486 ( .A0(n2355), .A1(n2371), .B0(n2354), .Y(n2373) );
  OR2X4 U1488 ( .A(n1095), .B(n1023), .Y(n1022) );
  CLKINVX3 U1489 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_2[4] ), .Y(n1023) );
  NAND2X4 U1490 ( .A(n2174), .B(n2177), .Y(n2168) );
  NAND2X6 U1491 ( .A(n2378), .B(n2377), .Y(n2400) );
  NAND2BX4 U1492 ( .AN(n2635), .B(n2634), .Y(n2637) );
  AND2X8 U1494 ( .A(n1010), .B(n798), .Y(n2338) );
  OAI21X2 U1495 ( .A0(n2633), .A1(n2632), .B0(n2631), .Y(n2634) );
  AOI21X8 U1496 ( .A0(n2589), .A1(n1235), .B0(n2598), .Y(n2603) );
  OAI2BB1X4 U1497 ( .A0N(n2423), .A1N(n2542), .B0(n2539), .Y(n2426) );
  XNOR2X4 U1499 ( .A(n2606), .B(n796), .Y(n2620) );
  OAI2B11X2 U1500 ( .A1N(n685), .A0(\decoder/w_PM_1[1] ), .B0(
        \decoder/w_PM_1[0] ), .C0(n1051), .Y(n2812) );
  MXI2X4 U1501 ( .A(n1563), .B(n1561), .S0(n1434), .Y(n669) );
  BUFX6 U1502 ( .A(n2172), .Y(n1122) );
  INVX2 U1503 ( .A(n683), .Y(n2823) );
  INVX2 U1505 ( .A(n1156), .Y(n1157) );
  AOI21X1 U1506 ( .A0(n709), .A1(n2808), .B0(n2803), .Y(n2816) );
  NAND2BX2 U1507 ( .AN(n2305), .B(n2306), .Y(n2232) );
  AOI21X1 U1508 ( .A0(n2840), .A1(n2839), .B0(n2838), .Y(n2841) );
  AOI31X1 U1509 ( .A0(n2898), .A1(n709), .A2(n2897), .B0(n2896), .Y(n2899) );
  INVX2 U1514 ( .A(n2238), .Y(n2217) );
  NAND2BX2 U1516 ( .AN(n1864), .B(n1863), .Y(n1867) );
  NAND2X4 U1517 ( .A(n2556), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[1] ), .Y(
        n2555) );
  NAND3X2 U1518 ( .A(n2545), .B(n1122), .C(n2171), .Y(n2173) );
  NAND2X4 U1520 ( .A(n1159), .B(n1160), .Y(n1161) );
  OAI2BB1X1 U1523 ( .A0N(n1462), .A1N(n1145), .B0(n2984), .Y(
        \decoder/u_cmp_sel/N42 ) );
  INVX6 U1526 ( .A(n2337), .Y(n2345) );
  OAI21X1 U1527 ( .A0(n1121), .A1(\decoder/w_PM_1[1] ), .B0(
        \decoder/w_PM_1[0] ), .Y(n1025) );
  NOR2XL U1528 ( .A(n699), .B(n1025), .Y(n2844) );
  OAI21X1 U1529 ( .A0(n2906), .A1(\decoder/w_PM_1[6] ), .B0(n2855), .Y(n1026)
         );
  AOI2B1X1 U1530 ( .A1N(n2850), .A0(n2827), .B0(n1026), .Y(n2801) );
  NOR2BX1 U1531 ( .AN(\decoder/u_ACS_matrix/w_PM_2_to_3_1[0] ), .B(
        \decoder/u_ACS_matrix/w_PM_2_to_3_2[0] ), .Y(n1761) );
  NAND4BX2 U1533 ( .AN(n2065), .B(n2066), .C(n2068), .D(n2996), .Y(n2069) );
  AND2X1 U1536 ( .A(n1664), .B(n1669), .Y(n1665) );
  INVX2 U1537 ( .A(n1620), .Y(n1028) );
  AOI2BB2XL U1538 ( .B0(n2142), .B1(n1042), .A0N(n1028), .A1N(n2141), .Y(n775)
         );
  AOI22XL U1539 ( .A0(n1616), .A1(\decoder/u_input_shifter/w_data_6[6] ), .B0(
        n2389), .B1(\decoder/u_input_shifter/w_data_1[6] ), .Y(n1029) );
  AOI22XL U1540 ( .A0(n1615), .A1(\decoder/u_input_shifter/w_data_4[6] ), .B0(
        n1614), .B1(\decoder/u_input_shifter/w_data_3[6] ), .Y(n1030) );
  AOI22XL U1541 ( .A0(n1617), .A1(\decoder/u_input_shifter/w_data_8[6] ), .B0(
        n2393), .B1(\decoder/u_input_shifter/w_data_7[6] ), .Y(n1031) );
  AOI22XL U1542 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_5[6] ), .B0(
        n1619), .B1(\decoder/u_input_shifter/w_data_2[6] ), .Y(n1032) );
  NAND4X2 U1543 ( .A(n1029), .B(n1030), .C(n1031), .D(n1032), .Y(
        \decoder/u_input_shifter/U_input_split/N43 ) );
  NAND2X2 U1544 ( .A(n1438), .B(n1440), .Y(n1033) );
  MXI2X4 U1545 ( .A(n1538), .B(n1536), .S0(n1033), .Y(n670) );
  OAI22X1 U1546 ( .A0(n1098), .A1(n698), .B0(n697), .B1(n2824), .Y(n1034) );
  NOR2X1 U1547 ( .A(n2826), .B(n1034), .Y(n1035) );
  OAI22X1 U1548 ( .A0(n685), .A1(n1121), .B0(n686), .B1(n2864), .Y(n1036) );
  NAND2X2 U1549 ( .A(n1035), .B(n1036), .Y(n2853) );
  OA21X2 U1552 ( .A0(\decoder/u_ACS_matrix/w_PM_3_to_4_4[0] ), .A1(n1804), 
        .B0(n1862), .Y(n1874) );
  NAND2XL U1554 ( .A(n2680), .B(n2681), .Y(n1038) );
  OAI21X1 U1555 ( .A0(n1038), .A1(n2683), .B0(n1037), .Y(n2685) );
  NAND2XL U1556 ( .A(n1757), .B(n1785), .Y(n1039) );
  INVXL U1557 ( .A(n863), .Y(n1040) );
  AOI31X1 U1558 ( .A0(n2042), .A1(n1040), .A2(n2050), .B0(n1937), .Y(n1983) );
  OAI2BB1X4 U1560 ( .A0N(n1894), .A1N(n1895), .B0(n1896), .Y(n1902) );
  AOI2BB1X2 U1561 ( .A0N(n1702), .A1N(n1164), .B0(n1665), .Y(n1671) );
  AOI21X2 U1562 ( .A0(n1693), .A1(n1696), .B0(n1692), .Y(n1041) );
  OA21X4 U1563 ( .A0(n1186), .A1(n1041), .B0(n1698), .Y(n1699) );
  INVX2 U1564 ( .A(n1620), .Y(n1042) );
  AOI22XL U1566 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_1[15] ), 
        .B0(n2389), .B1(\decoder/u_input_shifter/w_data_5[15] ), .Y(n1043) );
  AOI22XL U1567 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_7[15] ), 
        .B0(n2393), .B1(\decoder/u_input_shifter/w_data_3[15] ), .Y(n1044) );
  AOI22XL U1568 ( .A0(n1617), .A1(\decoder/u_input_shifter/w_data_4[15] ), 
        .B0(n1615), .B1(\decoder/u_input_shifter/w_data_8[15] ), .Y(n1045) );
  AOI22XL U1569 ( .A0(n1616), .A1(\decoder/u_input_shifter/w_data_2[15] ), 
        .B0(n1619), .B1(\decoder/u_input_shifter/w_data_6[15] ), .Y(n1046) );
  AND4X2 U1570 ( .A(n1043), .B(n1044), .C(n1045), .D(n1046), .Y(n342) );
  NOR2BX8 U1571 ( .AN(n324), .B(\decoder/w_enc_bit_3[0] ), .Y(n1708) );
  NAND2XL U1572 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_3[3] ), .B(
        \decoder/u_ACS_matrix/w_PM_6_to_7_3[2] ), .Y(n1047) );
  MXI2X1 U1573 ( .A(n2547), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[4] ), .S0(
        n1047), .Y(n2201) );
  NOR3X1 U1575 ( .A(n2167), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_4[3] ), .C(
        n2175), .Y(n1131) );
  NOR3BX1 U1576 ( .AN(\decoder/u_ACS_matrix/w_PM_7_to_8_3[2] ), .B(n2678), .C(
        n2715), .Y(n1048) );
  INVX2 U1578 ( .A(n1049), .Y(n1920) );
  OAI2B1X1 U1579 ( .A1N(n1667), .A0(\decoder/u_ACS_matrix/w_PM_1_to_2_1[0] ), 
        .B0(n1668), .Y(n1702) );
  INVXL U1581 ( .A(n1681), .Y(n1050) );
  AOI2BB2XL U1582 ( .B0(n1661), .B1(n1050), .A0N(n1050), .A1N(n1660), .Y(n931)
         );
  INVXL U1583 ( .A(n686), .Y(n1051) );
  NAND2BX1 U1584 ( .AN(n1772), .B(n1773), .Y(n1775) );
  CLKNAND2X2 U1586 ( .A(n2028), .B(n2083), .Y(n1052) );
  OAI2B11X2 U1588 ( .A1N(n2085), .A0(n2084), .B0(n1053), .C0(n1052), .Y(n2034)
         );
  INVXL U1591 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_4[5] ), .Y(n1055) );
  NAND3BXL U1595 ( .AN(n2505), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_2[4] ), 
        .C(n2438), .Y(n1057) );
  XOR2X1 U1596 ( .A(n2478), .B(n1057), .Y(n2519) );
  NOR2XL U1597 ( .A(n1216), .B(n1219), .Y(n1058) );
  NAND3X2 U1598 ( .A(n1218), .B(n1058), .C(n1217), .Y(n2749) );
  NAND3XL U1599 ( .A(n1993), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_4[3] ), .C(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[4] ), .Y(n1988) );
  OAI2B1X2 U1600 ( .A1N(n1702), .A0(n1188), .B0(n1704), .Y(n1705) );
  AND2X6 U1601 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_3[2] ), .B(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[1] ), .Y(n2723) );
  AOI2BB2XL U1604 ( .B0(n1620), .B1(n2144), .A0N(n2143), .A1N(n1620), .Y(n774)
         );
  AOI22XL U1605 ( .A0(n1615), .A1(\decoder/u_input_shifter/w_data_4[7] ), .B0(
        n1617), .B1(\decoder/u_input_shifter/w_data_8[7] ), .Y(n1059) );
  AOI22XL U1606 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_5[7] ), .B0(
        n1619), .B1(\decoder/u_input_shifter/w_data_2[7] ), .Y(n1060) );
  AOI22XL U1607 ( .A0(n1616), .A1(\decoder/u_input_shifter/w_data_6[7] ), .B0(
        n2389), .B1(\decoder/u_input_shifter/w_data_1[7] ), .Y(n1061) );
  AOI22XL U1608 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_3[7] ), .B0(
        n2393), .B1(\decoder/u_input_shifter/w_data_7[7] ), .Y(n1062) );
  AND4X2 U1609 ( .A(n1059), .B(n1060), .C(n1061), .D(n1062), .Y(n326) );
  NOR2BX1 U1610 ( .AN(n1698), .B(n1186), .Y(n938) );
  NOR3X1 U1613 ( .A(n2203), .B(n2201), .C(n1063), .Y(n2204) );
  NOR2BX1 U1615 ( .AN(n1763), .B(n1754), .Y(n1781) );
  CLKNAND2X2 U1616 ( .A(n1779), .B(n1778), .Y(n1791) );
  NAND2BX1 U1617 ( .AN(n2086), .B(n1859), .Y(n1320) );
  OAI2B1X1 U1618 ( .A1N(n2211), .A0(\decoder/u_ACS_matrix/w_PM_5_to_6_4[0] ), 
        .B0(n2219), .Y(n2311) );
  AOI2B1X1 U1619 ( .A1N(\decoder/u_ACS_matrix/w_PM_5_to_6_4[3] ), .A0(n2241), 
        .B0(n2242), .Y(n2303) );
  NOR2BX1 U1620 ( .AN(\decoder/u_ACS_matrix/w_PM_6_to_7_4[5] ), .B(n2207), .Y(
        n2376) );
  OAI2B1X1 U1621 ( .A1N(n1713), .A0(\decoder/u_ACS_matrix/w_PM_2_to_3_1[0] ), 
        .B0(n1752), .Y(n1787) );
  NOR2BX1 U1622 ( .AN(n732), .B(n1624), .Y(n705) );
  NAND3XL U1628 ( .A(n2737), .B(n2736), .C(n2713), .Y(n1065) );
  CLKNAND2X2 U1629 ( .A(n1065), .B(n2678), .Y(n2708) );
  AOI2B1X1 U1630 ( .A1N(n2326), .A0(n2328), .B0(n2215), .Y(n794) );
  OAI21X1 U1631 ( .A0(n1915), .A1(n982), .B0(n1914), .Y(n1066) );
  OAI21X1 U1632 ( .A0(n1917), .A1(n1132), .B0(n1066), .Y(n872) );
  AOI22XL U1633 ( .A0(n1616), .A1(\decoder/u_input_shifter/w_data_8[2] ), .B0(
        n2389), .B1(\decoder/u_input_shifter/w_data_3[2] ), .Y(n1067) );
  AOI22XL U1634 ( .A0(n1615), .A1(\decoder/u_input_shifter/w_data_6[2] ), .B0(
        n1614), .B1(\decoder/u_input_shifter/w_data_5[2] ), .Y(n1068) );
  AOI22XL U1635 ( .A0(n1617), .A1(\decoder/u_input_shifter/w_data_2[2] ), .B0(
        n2393), .B1(\decoder/u_input_shifter/w_data_1[2] ), .Y(n1069) );
  AOI22XL U1636 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_7[2] ), .B0(
        n1619), .B1(\decoder/u_input_shifter/w_data_4[2] ), .Y(n1070) );
  NAND4X1 U1637 ( .A(n1067), .B(n1068), .C(n1069), .D(n1070), .Y(
        \decoder/u_input_shifter/U_input_split/N39 ) );
  AND2X2 U1639 ( .A(n1436), .B(n1033), .Y(n1071) );
  INVXL U1640 ( .A(n1975), .Y(n2087) );
  INVXL U1642 ( .A(n1907), .Y(n1906) );
  MXI2X2 U1644 ( .A(n1470), .B(n1468), .S0(n1100), .Y(n683) );
  INVX4 U1645 ( .A(\decoder/u_ACS_matrix/w_PM_4_to_5_3[2] ), .Y(n1133) );
  INVXL U1646 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_3[1] ), .Y(n1738) );
  AND2X2 U1647 ( .A(n1315), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[2] ), .Y(
        n1074) );
  NAND2BX4 U1648 ( .AN(n2267), .B(n2258), .Y(n2320) );
  CLKBUFX4 U1650 ( .A(n3039), .Y(n1634) );
  INVX2 U1654 ( .A(n1080), .Y(n1272) );
  MXI2X2 U1656 ( .A(n1332), .B(n1330), .S0(n1082), .Y(n748) );
  INVXL U1661 ( .A(n1090), .Y(\decoder/u_ACS_matrix/w_PM_1_to_2_1[0] ) );
  INVX2 U1662 ( .A(n1090), .Y(\decoder/u_ACS_matrix/w_PM_1_to_2_3[0] ) );
  MXI2X6 U1669 ( .A(n1480), .B(n1478), .S0(n1476), .Y(n725) );
  INVX4 U1671 ( .A(n796), .Y(n1095) );
  MX2X4 U1675 ( .A(n1396), .B(n1394), .S0(n1100), .Y(n1098) );
  MXI2X4 U1676 ( .A(n1363), .B(n1361), .S0(n1100), .Y(n682) );
  CLKINVX3 U1677 ( .A(n681), .Y(n2799) );
  NAND2BXL U1678 ( .AN(\decoder/w_PM_2[5] ), .B(n681), .Y(n2850) );
  NAND2BXL U1679 ( .AN(n681), .B(\decoder/w_PM_2[5] ), .Y(n2828) );
  NAND2BX2 U1682 ( .AN(\decoder/u_ACS_matrix/w_PM_7_to_8_3[0] ), .B(n2737), 
        .Y(n1317) );
  NOR2X2 U1684 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_3[0] ), .B(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[2] ), .Y(n2719) );
  AOI2BB2X1 U1686 ( .B0(n2719), .B1(n2721), .A0N(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[2] ), .A1N(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[1] ), .Y(n1203) );
  INVX2 U1688 ( .A(n2706), .Y(n1103) );
  XNOR2X1 U1689 ( .A(n2678), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[2] ), .Y(
        n2706) );
  INVX2 U1690 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_3[2] ), .Y(n1202) );
  NAND2X2 U1691 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_3[4] ), .B(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[3] ), .Y(n2715) );
  INVX2 U1692 ( .A(n1177), .Y(n2645) );
  NAND2X2 U1695 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_2[0] ), .B(n2597), .Y(
        n2587) );
  XNOR2X4 U1696 ( .A(n1198), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_2[0] ), .Y(
        n2413) );
  OR2X4 U1698 ( .A(n1613), .B(n1248), .Y(n2225) );
  INVXL U1701 ( .A(\decoder/u_input_shifter/U_input_split/N51 ), .Y(n1108) );
  OAI2BB1X4 U1702 ( .A0N(\decoder/u_ACS_matrix/w_PM_7_to_8_2[0] ), .A1N(n1255), 
        .B0(n1210), .Y(n2431) );
  XNOR2X1 U1705 ( .A(\decoder/u_input_shifter/U_input_split/N49 ), .B(n338), 
        .Y(n1112) );
  NAND2BX2 U1706 ( .AN(n2178), .B(n1131), .Y(n2179) );
  CLKINVX1 U1712 ( .A(n2548), .Y(n1598) );
  NAND2X2 U1713 ( .A(n1117), .B(n1074), .Y(n2548) );
  CLKINVX1 U1714 ( .A(n2555), .Y(n1117) );
  NOR2X8 U1715 ( .A(n1145), .B(n2915), .Y(n2982) );
  NAND2BX8 U1716 ( .AN(n2913), .B(n2914), .Y(n1118) );
  OAI211X4 U1717 ( .A0(n1020), .A1(n2860), .B0(n2859), .C0(n2858), .Y(n2915)
         );
  BUFX4 U1718 ( .A(n748), .Y(n1144) );
  DLY1X1 U1719 ( .A(n1006), .Y(n1119) );
  NAND2BX8 U1720 ( .AN(n2170), .B(n2169), .Y(n2182) );
  NOR2X1 U1722 ( .A(n1793), .B(n1780), .Y(n920) );
  INVX4 U1724 ( .A(n1789), .Y(n1793) );
  INVX1 U1726 ( .A(n1791), .Y(n1792) );
  NOR2BX2 U1727 ( .AN(n1730), .B(n1764), .Y(n912) );
  NOR2X4 U1729 ( .A(n1238), .B(n2071), .Y(n2075) );
  INVX5 U1730 ( .A(n2079), .Y(n2940) );
  INVX6 U1731 ( .A(n1820), .Y(n2920) );
  OAI2BB1X2 U1732 ( .A0N(n2575), .A1N(n2569), .B0(n2572), .Y(n1276) );
  XNOR2X2 U1735 ( .A(n2507), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_1[5] ), .Y(
        n2531) );
  CLKINVX4 U1736 ( .A(n2289), .Y(n2288) );
  CLKINVX4 U1739 ( .A(n2475), .Y(n2507) );
  INVX2 U1740 ( .A(n2063), .Y(n2097) );
  INVXL U1741 ( .A(n1819), .Y(n1821) );
  INVX2 U1742 ( .A(n2196), .Y(n2381) );
  INVX4 U1743 ( .A(n958), .Y(n1152) );
  NAND2X4 U1744 ( .A(n2263), .B(n1157), .Y(n2276) );
  INVXL U1745 ( .A(n2683), .Y(n2671) );
  MXI2XL U1746 ( .A(n1188), .B(n1706), .S0(n1705), .Y(n942) );
  NOR2X1 U1747 ( .A(n1731), .B(n1747), .Y(n1748) );
  MXI2XL U1748 ( .A(n1703), .B(n1702), .S0(n1705), .Y(n943) );
  INVXL U1750 ( .A(n1794), .Y(n1796) );
  INVX1 U1753 ( .A(n1140), .Y(n1141) );
  INVX1 U1754 ( .A(n342), .Y(n1528) );
  INVXL U1755 ( .A(n1731), .Y(n1746) );
  NOR2X1 U1756 ( .A(n2065), .B(n2042), .Y(n1947) );
  INVX1 U1757 ( .A(n1719), .Y(n1716) );
  CLKNAND2X2 U1758 ( .A(\decoder/u_input_shifter/U_input_split/N51 ), .B(n342), 
        .Y(n1591) );
  INVX1 U1759 ( .A(n1146), .Y(n1147) );
  INVX1 U1760 ( .A(n1729), .Y(n1788) );
  NAND2X4 U1762 ( .A(n2345), .B(n796), .Y(n2346) );
  INVX1 U1763 ( .A(n2690), .Y(n2697) );
  NAND2X1 U1764 ( .A(n1660), .B(n1661), .Y(n1594) );
  INVXL U1765 ( .A(n1704), .Y(n1706) );
  CLKNAND2X2 U1766 ( .A(n1732), .B(n1865), .Y(n1733) );
  OAI2BB1XL U1767 ( .A0N(n1864), .A1N(n1874), .B0(n1883), .Y(n1740) );
  INVX1 U1768 ( .A(n2094), .Y(n2053) );
  CLKNAND2X2 U1769 ( .A(n1668), .B(n1664), .Y(n1704) );
  INVX1 U1770 ( .A(n1660), .Y(n1680) );
  INVXL U1773 ( .A(n1695), .Y(n1659) );
  NOR2X1 U1774 ( .A(n2551), .B(n1316), .Y(n2552) );
  INVX1 U1775 ( .A(n2866), .Y(n2867) );
  INVX1 U1776 ( .A(n1559), .Y(n2820) );
  CLKINVX4 U1778 ( .A(n1231), .Y(n1894) );
  NAND2X1 U1779 ( .A(n2260), .B(n2259), .Y(n2261) );
  CLKNAND2X2 U1780 ( .A(n2828), .B(n2827), .Y(n2849) );
  AO21X1 U1781 ( .A0(n465), .A1(n1640), .B0(
        \decoder/u_input_shifter/u_input_fifo/N28 ), .Y(n463) );
  NOR2XL U1782 ( .A(n2259), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[1] ), .Y(
        n2106) );
  INVX2 U1783 ( .A(n2558), .Y(n2580) );
  INVX1 U1785 ( .A(n2343), .Y(n2341) );
  AOI21XL U1786 ( .A0(n1643), .A1(n1644), .B0(n2389), .Y(n345) );
  NAND2X1 U1787 ( .A(n2030), .B(n2029), .Y(n2031) );
  CLKNAND2X2 U1788 ( .A(n2805), .B(n2804), .Y(n2803) );
  INVX1 U1789 ( .A(n2808), .Y(n2807) );
  NOR2X1 U1790 ( .A(n2029), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_1[1] ), .Y(
        n1844) );
  MXI2XL U1791 ( .A(n1424), .B(n1422), .S0(n2976), .Y(n718) );
  INVXL U1792 ( .A(n1168), .Y(n1215) );
  INVXL U1793 ( .A(n1166), .Y(n1212) );
  INVXL U1794 ( .A(n1169), .Y(n1214) );
  INVXL U1795 ( .A(n1167), .Y(n1213) );
  NOR2X1 U1796 ( .A(n1636), .B(n484), .Y(n950) );
  NOR2X1 U1797 ( .A(n1641), .B(n1639), .Y(
        \decoder/u_input_shifter/u_input_fifo/N8 ) );
  NOR2X1 U1798 ( .A(n1640), .B(n1639), .Y(n949) );
  NOR2X1 U1799 ( .A(n484), .B(n1638), .Y(n948) );
  NOR2X1 U1800 ( .A(n465), .B(n1641), .Y(n952) );
  NOR2X1 U1801 ( .A(n2023), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_1[1] ), .Y(
        n2026) );
  NAND2XL U1802 ( .A(n1640), .B(n1641), .Y(n482) );
  MXI2XL U1803 ( .A(n1371), .B(n1369), .S0(n2976), .Y(n716) );
  MXI2XL U1804 ( .A(n1375), .B(n1373), .S0(n2976), .Y(n715) );
  INVXL U1805 ( .A(n1696), .Y(n1658) );
  MXI2XL U1806 ( .A(n1379), .B(n1377), .S0(n2976), .Y(n714) );
  MXI2XL U1808 ( .A(n1367), .B(n1365), .S0(n2976), .Y(n717) );
  INVXL U1809 ( .A(n2985), .Y(
        \decoder/u_ACS_matrix/u_ACS_col_1/u_ACS_mem_3/u_ACS/ham_dist_2[0] ) );
  INVXL U1810 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_4[4] ), .Y(n1987) );
  INVX1 U1811 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_4[5] ), .Y(n2570) );
  INVXL U1812 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_3[4] ), .Y(n2717) );
  INVX1 U1813 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_3[2] ), .Y(n2971) );
  INVX1 U1814 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_4[2] ), .Y(n2970) );
  NAND2X2 U1815 ( .A(n484), .B(n487), .Y(n1641) );
  INVXL U1816 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_2[4] ), .Y(n2119) );
  INVX1 U1817 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_1[1] ), .Y(n1271) );
  INVXL U1819 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_1[4] ), .Y(n2436) );
  CLKNAND2X2 U1820 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_1[1] ), .B(
        \decoder/u_ACS_matrix/w_PM_5_to_6_1[2] ), .Y(n2265) );
  INVXL U1821 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_4[3] ), .Y(n1990) );
  INVX1 U1822 ( .A(\decoder/w_PM_1[0] ), .Y(n2886) );
  MXI2X4 U1823 ( .A(n1336), .B(n1334), .S0(n1102), .Y(n695) );
  INVXL U1824 ( .A(n484), .Y(n1637) );
  INVXL U1826 ( .A(\decoder/u_ACS_matrix/w_PM_2_to_3_4[1] ), .Y(n1768) );
  OR2X2 U1827 ( .A(n313), .B(\decoder/w_enc_bit_2[0] ), .Y(n1696) );
  INVX1 U1828 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_4[5] ), .Y(n2794) );
  INVX1 U1829 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_4[4] ), .Y(n2931) );
  INVX1 U1830 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_4[3] ), .Y(n2947) );
  INVX1 U1831 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_4[2] ), .Y(n2958) );
  INVX2 U1832 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_1[2] ), .Y(n2482) );
  INVX1 U1833 ( .A(\decoder/w_PM_2[5] ), .Y(n2835) );
  INVX1 U1834 ( .A(\decoder/w_PM_4[6] ), .Y(n2904) );
  INVXL U1835 ( .A(n1897), .Y(n1806) );
  INVX1 U1836 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_2[0] ), .Y(n1803) );
  NAND3X4 U1837 ( .A(n1263), .B(n1262), .C(n2196), .Y(n2206) );
  NAND3X4 U1838 ( .A(n1130), .B(n2187), .C(n2186), .Y(n1263) );
  NAND2X2 U1839 ( .A(n1123), .B(n2526), .Y(n2492) );
  NAND2X4 U1840 ( .A(n2532), .B(n2512), .Y(n2513) );
  OAI22X2 U1841 ( .A0(n2569), .A1(n2575), .B0(n2581), .B1(n1279), .Y(n1278) );
  AOI2BB2X2 U1842 ( .B0(n2486), .B1(n2429), .A0N(n2428), .A1N(n1271), .Y(n2528) );
  NAND2X4 U1844 ( .A(n1305), .B(n1243), .Y(n1304) );
  CLKNAND2X2 U1845 ( .A(n2541), .B(n2497), .Y(n2495) );
  NAND2X4 U1846 ( .A(n2619), .B(n2590), .Y(n2596) );
  NAND2X4 U1847 ( .A(n2431), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_2[1] ), .Y(
        n2430) );
  NOR2X6 U1850 ( .A(n2416), .B(n2415), .Y(n2448) );
  OAI21X2 U1851 ( .A0(n2438), .A1(\decoder/u_ACS_matrix/w_PM_7_to_8_2[4] ), 
        .B0(n2461), .Y(n2712) );
  NAND2X4 U1854 ( .A(n1237), .B(n1209), .Y(n1236) );
  NAND3X2 U1855 ( .A(n2446), .B(n2445), .C(n2455), .Y(n2457) );
  XNOR2X2 U1856 ( .A(n2451), .B(n2450), .Y(n2533) );
  NOR2X4 U1857 ( .A(n2196), .B(n2380), .Y(n1260) );
  OAI21X2 U1858 ( .A0(\decoder/u_ACS_matrix/w_PM_6_to_7_3[3] ), .A1(n2188), 
        .B0(n2190), .Y(n2383) );
  MXI2X4 U1860 ( .A(n1426), .B(n1428), .S0(n1272), .Y(n711) );
  AO2B2X4 U1861 ( .B0(n2890), .B1(n711), .A0(\decoder/w_PM_1[3] ), .A1N(n669), 
        .Y(n2893) );
  NAND2X4 U1862 ( .A(n2174), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_4[1] ), .Y(
        n1305) );
  NAND2X4 U1863 ( .A(n2732), .B(n2737), .Y(n2733) );
  NAND2X8 U1864 ( .A(n2338), .B(n797), .Y(n2337) );
  OAI2BB1X1 U1868 ( .A0N(n1128), .A1N(n2586), .B0(n2334), .Y(n2411) );
  INVXL U1869 ( .A(n1010), .Y(n1128) );
  NAND2X4 U1870 ( .A(n1304), .B(n2168), .Y(n1303) );
  NAND2X8 U1871 ( .A(n2597), .B(n2604), .Y(n2340) );
  OAI21X2 U1873 ( .A0(n2558), .A1(n2579), .B0(n1000), .Y(n1269) );
  NAND2X4 U1874 ( .A(n2564), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_4[3] ), .Y(
        n2563) );
  INVX6 U1875 ( .A(n2172), .Y(n2557) );
  NOR2X4 U1876 ( .A(n2384), .B(n1302), .Y(n2187) );
  NAND2BX8 U1879 ( .AN(n2178), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[0] ), 
        .Y(n2545) );
  OR2X4 U1880 ( .A(n1891), .B(n1894), .Y(n1892) );
  AO21X4 U1881 ( .A0(n1911), .A1(n1916), .B0(n1915), .Y(n1132) );
  NAND3X4 U1882 ( .A(n1226), .B(n1777), .C(n1225), .Y(n1779) );
  NOR2X8 U1883 ( .A(\decoder/w_enc_bit_5[0] ), .B(n332), .Y(n2066) );
  OAI2B1X4 U1886 ( .A1N(n1779), .A0(n1771), .B0(n1791), .Y(n1789) );
  OAI21X8 U1887 ( .A0(n1309), .A1(n2009), .B0(n1308), .Y(n1620) );
  AOI21X4 U1888 ( .A0(n2005), .A1(n2006), .B0(n2004), .Y(n1309) );
  NAND2BX4 U1889 ( .AN(n2239), .B(n2243), .Y(n2245) );
  OAI2BB1X4 U1894 ( .A0N(n1888), .A1N(n1887), .B0(n1886), .Y(n1924) );
  CLKINVX3 U1895 ( .A(n2721), .Y(n2724) );
  NAND2XL U1897 ( .A(n2141), .B(n2142), .Y(n2002) );
  NAND2X4 U1899 ( .A(n1782), .B(n1593), .Y(n1786) );
  AOI21X1 U1901 ( .A0(n2144), .A1(n2143), .B0(n2000), .Y(n2001) );
  OAI21X2 U1903 ( .A0(n1682), .A1(\decoder/u_ACS_matrix/w_PM_2_to_3_4[1] ), 
        .B0(n1687), .Y(n1725) );
  AOI31X4 U1904 ( .A0(n1718), .A1(n1717), .A2(n1259), .B0(n1192), .Y(n1730) );
  OAI2B2X2 U1905 ( .A1N(n1287), .A0(n1160), .B0(n2314), .B1(n2313), .Y(n807)
         );
  NOR2BX1 U1908 ( .AN(\decoder/u_ACS_matrix/w_data_5_to_6_4[1] ), .B(n2964), 
        .Y(n803) );
  INVX2 U1909 ( .A(n2023), .Y(n1135) );
  NOR2X2 U1910 ( .A(n2048), .B(n2047), .Y(n2052) );
  INVX4 U1912 ( .A(n2320), .Y(n1136) );
  CLKINVX3 U1913 ( .A(n1933), .Y(n1949) );
  NAND2X6 U1914 ( .A(n1934), .B(n861), .Y(n1933) );
  AOI21X6 U1916 ( .A0(n1264), .A1(n2255), .B0(n2256), .Y(n2267) );
  INVX6 U1918 ( .A(n798), .Y(n2586) );
  OAI21X1 U1919 ( .A0(n1934), .A1(n861), .B0(n1933), .Y(n1138) );
  OAI21X2 U1920 ( .A0(n1977), .A1(n1979), .B0(n1944), .Y(n1945) );
  OAI21X2 U1921 ( .A0(n2891), .A1(\decoder/w_PM_1[3] ), .B0(n2897), .Y(n2901)
         );
  NAND2X2 U1922 ( .A(n2643), .B(n2620), .Y(n2630) );
  INVXL U1923 ( .A(n1982), .Y(n1140) );
  NAND2BX2 U1930 ( .AN(n2907), .B(n2883), .Y(n2885) );
  NAND2BX4 U1932 ( .AN(n2485), .B(n1312), .Y(n1310) );
  NOR2X4 U1933 ( .A(n1209), .B(n2437), .Y(n2438) );
  INVX4 U1934 ( .A(n1236), .Y(n2423) );
  OAI21X2 U1936 ( .A0(n2221), .A1(\decoder/u_ACS_matrix/w_PM_5_to_6_4[2] ), 
        .B0(n2241), .Y(n2306) );
  NAND3X4 U1939 ( .A(n2501), .B(n2500), .C(n2499), .Y(n2504) );
  OAI22X1 U1940 ( .A0(n2864), .A1(n672), .B0(n1121), .B1(n671), .Y(n2865) );
  INVXL U1941 ( .A(n2703), .Y(n2705) );
  NOR2X2 U1943 ( .A(n1961), .B(n1959), .Y(n1840) );
  NAND2XL U1944 ( .A(n2081), .B(n2078), .Y(n2015) );
  NAND3X4 U1950 ( .A(n1689), .B(n1688), .C(n1690), .Y(n1723) );
  BUFX6 U1951 ( .A(n2287), .Y(n1241) );
  INVXL U1953 ( .A(n1024), .Y(n1146) );
  NAND3X2 U1954 ( .A(n2108), .B(n2262), .C(n2107), .Y(n2111) );
  NAND2X4 U1955 ( .A(n2116), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_2[1] ), .Y(
        n2103) );
  NOR2BX4 U1957 ( .AN(n2424), .B(n2448), .Y(n2537) );
  NAND2BX2 U1958 ( .AN(\decoder/u_ACS_matrix/w_PM_7_to_8_1[3] ), .B(n2416), 
        .Y(n2424) );
  NAND2X4 U1960 ( .A(n2224), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_3[1] ), .Y(
        n2223) );
  OAI2B11X2 U1961 ( .A1N(n2578), .A0(n2577), .B0(n2562), .C0(n2561), .Y(n2568)
         );
  INVXL U1962 ( .A(n2745), .Y(n2782) );
  OAI21X2 U1963 ( .A0(n1713), .A1(\decoder/u_ACS_matrix/w_PM_2_to_3_3[0] ), 
        .B0(n1766), .Y(n1797) );
  NAND2BX8 U1964 ( .AN(n2211), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_4[0] ), 
        .Y(n2219) );
  XNOR2X4 U1966 ( .A(n2449), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_1[6] ), .Y(
        n2518) );
  INVX4 U1969 ( .A(n748), .Y(n2437) );
  INVX2 U1971 ( .A(n2057), .Y(n2058) );
  MXI2X6 U1972 ( .A(n1577), .B(n1575), .S0(n1573), .Y(n726) );
  XNOR2X4 U1974 ( .A(n2571), .B(n2570), .Y(n2573) );
  NAND2X4 U1975 ( .A(n2267), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_2[2] ), .Y(
        n2287) );
  OAI21X2 U1976 ( .A0(\decoder/u_ACS_matrix/w_PM_5_to_6_2[2] ), .A1(n2267), 
        .B0(n2287), .Y(n2318) );
  XNOR2X4 U1977 ( .A(n2287), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_2[3] ), .Y(
        n2315) );
  XNOR2X4 U1979 ( .A(n2677), .B(n2752), .Y(n2702) );
  OAI2BB1X4 U1980 ( .A0N(\decoder/w_enc_bit_8[0] ), .A1N(n1211), .B0(n1609), 
        .Y(n1210) );
  INVX2 U1981 ( .A(n2423), .Y(n2543) );
  AOI22X2 U1982 ( .A0(n2982), .A1(n701), .B0(n1145), .B1(\decoder/w_data_4[6] ), .Y(n2935) );
  AOI22X2 U1983 ( .A0(n2982), .A1(n703), .B0(\decoder/w_data_4[4] ), .B1(n1145), .Y(n2963) );
  AOI22X2 U1984 ( .A0(n2982), .A1(n702), .B0(\decoder/w_data_4[5] ), .B1(n1145), .Y(n2951) );
  OAI2B11X2 U1988 ( .A1N(n1975), .A0(n1860), .B0(n1319), .C0(n1321), .Y(n833)
         );
  NAND3X4 U1989 ( .A(n1857), .B(n1856), .C(n1858), .Y(n1860) );
  NAND2BX2 U1990 ( .AN(n1320), .B(n1860), .Y(n1319) );
  NAND2BX4 U1991 ( .AN(n1292), .B(n1291), .Y(n1624) );
  XNOR2X4 U1992 ( .A(n2419), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_1[2] ), .Y(
        n2542) );
  INVX4 U1993 ( .A(n2195), .Y(n2380) );
  NOR2XL U1994 ( .A(n2375), .B(n2195), .Y(n2193) );
  XNOR2X4 U1995 ( .A(n2207), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_4[5] ), .Y(
        n2195) );
  NAND2X8 U1997 ( .A(n1893), .B(n1897), .Y(n1804) );
  AND3X6 U1998 ( .A(n2180), .B(n2179), .C(n1294), .Y(n2384) );
  NAND3X2 U1999 ( .A(n2853), .B(n2852), .C(n2829), .Y(n2830) );
  OAI211X4 U2000 ( .A0(n2816), .A1(n2815), .B0(n2814), .C0(n2813), .Y(n2832)
         );
  INVX2 U2001 ( .A(n2059), .Y(n1154) );
  OAI21X4 U2002 ( .A0(n797), .A1(n2338), .B0(n2337), .Y(n2409) );
  NOR2X4 U2003 ( .A(n2555), .B(n2549), .Y(n2566) );
  AOI2BB2X4 U2004 ( .B0(n2877), .B1(n2876), .A0N(n2875), .A1N(n2874), .Y(n2914) );
  OAI21X2 U2005 ( .A0(n2554), .A1(\decoder/u_ACS_matrix/w_PM_6_to_7_4[1] ), 
        .B0(n2553), .Y(n2578) );
  OAI21X2 U2006 ( .A0(\decoder/u_ACS_matrix/w_PM_4_to_5_3[1] ), .A1(n1939), 
        .B0(n1938), .Y(n1984) );
  NAND2X4 U2007 ( .A(n1939), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_3[1] ), .Y(
        n1938) );
  NAND3X8 U2008 ( .A(n1227), .B(n2246), .C(n2247), .Y(n2964) );
  NAND3X4 U2009 ( .A(n1230), .B(n2245), .C(n2304), .Y(n2246) );
  NOR2X4 U2010 ( .A(n2223), .B(n2218), .Y(n2238) );
  NAND2X4 U2011 ( .A(n1196), .B(n2349), .Y(n2405) );
  NAND2X4 U2012 ( .A(n2642), .B(n2596), .Y(n2612) );
  CLKINVX3 U2014 ( .A(n2783), .Y(n2766) );
  NAND3X4 U2017 ( .A(n2771), .B(n2770), .C(n2775), .Y(n2777) );
  NAND3X2 U2018 ( .A(n1202), .B(n3067), .C(n2721), .Y(n1201) );
  XNOR2X4 U2020 ( .A(n2127), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[4] ), .Y(
        n2151) );
  NAND3X4 U2021 ( .A(n2463), .B(n2462), .C(n2519), .Y(n2523) );
  NAND2X4 U2023 ( .A(n1999), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_3[1] ), .Y(
        n1998) );
  XNOR2X4 U2024 ( .A(n2007), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_3[4] ), .Y(
        n2162) );
  XNOR2X4 U2026 ( .A(n1843), .B(n1842), .Y(n1966) );
  NAND2X2 U2029 ( .A(n2262), .B(n2261), .Y(n1156) );
  NAND2X4 U2030 ( .A(n2297), .B(n2314), .Y(n1158) );
  NAND2BX4 U2031 ( .AN(n2322), .B(n2323), .Y(n2262) );
  AOI31X2 U2032 ( .A0(n2276), .A1(n2268), .A2(n2319), .B0(n1018), .Y(n2283) );
  NAND2X4 U2033 ( .A(n2325), .B(n2324), .Y(n2314) );
  NAND3X4 U2035 ( .A(n2296), .B(n2312), .C(n2295), .Y(n2297) );
  NAND2X4 U2037 ( .A(n1932), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_3[0] ), .Y(
        n2043) );
  XNOR2X4 U2039 ( .A(n2448), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_1[4] ), .Y(
        n2711) );
  AOI21X2 U2041 ( .A0(n1948), .A1(n1943), .B0(n1942), .Y(n1944) );
  OAI21X2 U2042 ( .A0(n2556), .A1(\decoder/u_ACS_matrix/w_PM_6_to_7_3[1] ), 
        .B0(n2555), .Y(n2577) );
  NAND2X4 U2043 ( .A(n1860), .B(n1859), .Y(n1956) );
  NOR2BX4 U2044 ( .AN(n2335), .B(n2333), .Y(n2342) );
  NAND2X2 U2045 ( .A(n2331), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_1[1] ), .Y(
        n2335) );
  NAND3X4 U2047 ( .A(n2469), .B(n2470), .C(n2518), .Y(n2522) );
  NAND2X4 U2048 ( .A(n1770), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_3[1] ), .Y(
        n1771) );
  INVX4 U2049 ( .A(n2296), .Y(n1159) );
  NAND3X4 U2052 ( .A(n1265), .B(n1266), .C(n2375), .Y(n2377) );
  MXI2X2 U2053 ( .A(n1519), .B(n1517), .S0(n1434), .Y(n668) );
  AOI21X4 U2055 ( .A0(n2073), .A1(n2072), .B0(n2062), .Y(n1238) );
  NOR2XL U2056 ( .A(n2488), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_1[1] ), .Y(
        n2429) );
  OAI21X8 U2057 ( .A0(n1933), .A1(n1955), .B0(n1976), .Y(n2952) );
  XNOR2X4 U2058 ( .A(n1142), .B(n1247), .Y(n2647) );
  NOR2X4 U2059 ( .A(\decoder/w_enc_bit_7[0] ), .B(n1611), .Y(n2546) );
  XNOR2X4 U2060 ( .A(n2190), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[4] ), .Y(
        n2196) );
  NAND2BX4 U2063 ( .AN(n2901), .B(n2893), .Y(n2900) );
  NAND2X4 U2064 ( .A(n2074), .B(n2097), .Y(n2098) );
  NAND3X2 U2065 ( .A(n2257), .B(n2256), .C(n1314), .Y(n2258) );
  NAND2BX4 U2066 ( .AN(n2536), .B(n2535), .Y(n2500) );
  NOR2X2 U2067 ( .A(n709), .B(n2845), .Y(n2837) );
  NAND4BXL U2068 ( .AN(n709), .B(n2805), .C(n682), .D(n2804), .Y(n2800) );
  MXI2X4 U2069 ( .A(n1484), .B(n1482), .S0(n1080), .Y(n709) );
  DLY1X1 U2070 ( .A(n3005), .Y(n1232) );
  NAND3X4 U2071 ( .A(n2060), .B(n2064), .C(n2068), .Y(n2073) );
  NAND2BX4 U2072 ( .AN(n2057), .B(n861), .Y(n2063) );
  OAI2BB1X2 U2073 ( .A0N(n1984), .A1N(n1983), .B0(n2051), .Y(n1943) );
  XNOR2X4 U2075 ( .A(n2603), .B(n2602), .Y(n1177) );
  NAND3X2 U2077 ( .A(n2269), .B(n2315), .C(n2276), .Y(n2280) );
  NOR2X2 U2078 ( .A(n3035), .B(n2318), .Y(n2269) );
  NAND3X4 U2079 ( .A(n2510), .B(n2509), .C(n2508), .Y(n2515) );
  NAND3X4 U2080 ( .A(n2504), .B(n2503), .C(n2502), .Y(n2510) );
  AOI21X2 U2082 ( .A0(n1982), .A1(n1980), .B0(n1940), .Y(n1948) );
  MXI2X6 U2083 ( .A(n1544), .B(n1542), .S0(n1433), .Y(n671) );
  OAI211X2 U2084 ( .A0(n1875), .A1(n1869), .B0(n1885), .C0(n1884), .Y(n1886)
         );
  NAND3X2 U2085 ( .A(n2277), .B(n2276), .C(n2315), .Y(n2278) );
  NOR2X2 U2086 ( .A(n3035), .B(n2274), .Y(n2277) );
  NAND3X4 U2088 ( .A(n3025), .B(n2255), .C(
        \decoder/u_ACS_matrix/w_PM_5_to_6_2[0] ), .Y(n2257) );
  NOR2X2 U2089 ( .A(n2823), .B(n669), .Y(n1559) );
  MXI2X6 U2090 ( .A(n1492), .B(n1490), .S0(n1100), .Y(n681) );
  INVX2 U2091 ( .A(n2275), .Y(n2268) );
  INVX2 U2093 ( .A(n2307), .Y(n2309) );
  CLKBUFX4 U2094 ( .A(n2395), .Y(n1618) );
  NAND2X2 U2096 ( .A(n1707), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_1[0] ), .Y(
        n1752) );
  INVX2 U2097 ( .A(n2773), .Y(n2774) );
  NOR2X2 U2102 ( .A(n1300), .B(n1298), .Y(n2727) );
  NOR2XL U2103 ( .A(n2952), .B(n1173), .Y(n825) );
  INVX2 U2105 ( .A(n2691), .Y(n2694) );
  NOR2BX1 U2106 ( .AN(n732), .B(n3092), .Y(n692) );
  INVX2 U2107 ( .A(n2583), .Y(n2584) );
  NAND2X2 U2108 ( .A(n1279), .B(n2581), .Y(n2567) );
  AOI21X2 U2110 ( .A0(\decoder/u_ACS_matrix/w_PM_6_to_7_4[0] ), .A1(n2340), 
        .B0(n2557), .Y(n2551) );
  OAI2BB1X2 U2112 ( .A0N(n2528), .A1N(n2530), .B0(n2434), .Y(n2445) );
  INVX2 U2115 ( .A(n2168), .Y(n1250) );
  INVX2 U2116 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_4[2] ), .Y(n1243) );
  AO22X2 U2117 ( .A0(n1076), .A1(n1581), .B0(n1579), .B1(n1088), .Y(n890) );
  NAND2X2 U2118 ( .A(n1800), .B(n1812), .Y(n1816) );
  INVX2 U2119 ( .A(n1812), .Y(n1817) );
  INVX2 U2120 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_2[2] ), .Y(n1908) );
  NOR2XL U2121 ( .A(n2351), .B(n2404), .Y(n2352) );
  NAND2BX2 U2122 ( .AN(n2117), .B(n2116), .Y(n2121) );
  NAND4X2 U2123 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_2[2] ), .B(
        \decoder/u_ACS_matrix/w_PM_5_to_6_2[1] ), .C(
        \decoder/u_ACS_matrix/w_PM_5_to_6_2[4] ), .D(
        \decoder/u_ACS_matrix/w_PM_5_to_6_2[3] ), .Y(n2117) );
  OAI21X1 U2124 ( .A0(\decoder/w_PM_4[6] ), .A1(n2872), .B0(n2871), .Y(n2880)
         );
  NAND2BX2 U2125 ( .AN(n667), .B(\decoder/w_PM_2[5] ), .Y(n2871) );
  INVX2 U2126 ( .A(\decoder/w_PM_1[1] ), .Y(n2887) );
  CLKINVX3 U2129 ( .A(n2485), .Y(n1311) );
  NAND2X4 U2130 ( .A(n2474), .B(n956), .Y(n2485) );
  INVX2 U2133 ( .A(n1952), .Y(n1955) );
  NOR2X2 U2134 ( .A(n2271), .B(n2270), .Y(n2272) );
  NOR2X2 U2135 ( .A(n2318), .B(n2274), .Y(n2273) );
  INVXL U2136 ( .A(n3025), .Y(n2250) );
  NAND2X2 U2137 ( .A(n2630), .B(n2629), .Y(n2623) );
  NOR2X2 U2138 ( .A(n2616), .B(n3096), .Y(n2633) );
  NOR2X2 U2139 ( .A(n2605), .B(n1155), .Y(n2610) );
  NAND3X2 U2141 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_1[0] ), .B(n2597), .C(
        n2604), .Y(n2599) );
  INVXL U2142 ( .A(n1983), .Y(n1985) );
  INVXL U2144 ( .A(n1980), .Y(n1981) );
  INVXL U2145 ( .A(n2692), .Y(n2693) );
  NAND3X4 U2147 ( .A(n1268), .B(n1267), .C(n2376), .Y(n2378) );
  AO22X4 U2150 ( .A0(n1076), .A1(n1585), .B0(n1583), .B1(n1088), .Y(n891) );
  NOR2BX4 U2151 ( .AN(\decoder/u_ACS_matrix/w_PM_3_to_4_2[0] ), .B(n1804), .Y(
        n1891) );
  OAI211X2 U2153 ( .A0(n2890), .A1(n711), .B0(n2889), .C0(n2888), .Y(n2902) );
  OAI2BB1X2 U2154 ( .A0N(n2487), .A1N(n2486), .B0(n2485), .Y(n2526) );
  NAND3X4 U2155 ( .A(n1311), .B(n1312), .C(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[4] ), .Y(n2475) );
  NOR2BX4 U2156 ( .AN(\decoder/u_ACS_matrix/w_PM_7_to_8_1[3] ), .B(n2482), .Y(
        n1312) );
  NAND3X4 U2157 ( .A(n2473), .B(n2432), .C(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[0] ), .Y(n2486) );
  NOR2BX2 U2158 ( .AN(n2089), .B(n2088), .Y(n2065) );
  MXI2X4 U2159 ( .A(n1349), .B(n1347), .S0(n978), .Y(n861) );
  CLKINVX3 U2160 ( .A(n1936), .Y(n1934) );
  NAND2X4 U2161 ( .A(n2254), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_2[0] ), .Y(
        n1264) );
  INVXL U2163 ( .A(n1964), .Y(n1965) );
  INVXL U2164 ( .A(n2528), .Y(n2529) );
  NAND3X2 U2165 ( .A(n2672), .B(n2703), .C(n2671), .Y(n2675) );
  OR2X4 U2168 ( .A(n2349), .B(n2594), .Y(n2401) );
  INVX2 U2171 ( .A(n709), .Y(n2878) );
  INVX2 U2172 ( .A(n2531), .Y(n2512) );
  XNOR2X4 U2174 ( .A(n2476), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_1[6] ), .Y(
        n2521) );
  NAND2X4 U2175 ( .A(n1954), .B(n1953), .Y(n1976) );
  INVXL U2176 ( .A(n2255), .Y(n2259) );
  OAI21X2 U2177 ( .A0(n2211), .A1(\decoder/u_ACS_matrix/w_PM_5_to_6_1[0] ), 
        .B0(n2252), .Y(n2323) );
  INVX2 U2179 ( .A(n2591), .Y(n2619) );
  XNOR2X4 U2180 ( .A(n1297), .B(n2593), .Y(n2656) );
  AND2X6 U2181 ( .A(n2603), .B(n1296), .Y(n2591) );
  MXI2X6 U2182 ( .A(n1342), .B(n1340), .S0(n1338), .Y(n798) );
  BUFX2 U2183 ( .A(n2388), .Y(n1616) );
  BUFX2 U2184 ( .A(n2390), .Y(n1615) );
  INVXL U2185 ( .A(n2699), .Y(n2701) );
  INVXL U2187 ( .A(n2569), .Y(n2576) );
  OAI21BX4 U2188 ( .A0(n1277), .A1(n1276), .B0N(n1275), .Y(n1293) );
  NAND2XL U2189 ( .A(n2583), .B(n2585), .Y(n2561) );
  NAND2X2 U2192 ( .A(n2432), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_2[0] ), .Y(
        n1256) );
  INVXL U2193 ( .A(n2379), .Y(n2208) );
  NAND3X2 U2194 ( .A(n1244), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_4[3] ), .C(
        n2181), .Y(n2180) );
  NAND2XL U2195 ( .A(n2983), .B(\decoder/w_data_3[5] ), .Y(n2950) );
  NAND2XL U2196 ( .A(n2983), .B(\decoder/w_data_3[4] ), .Y(n2962) );
  OAI211X2 U2197 ( .A0(n2360), .A1(n2361), .B0(n2359), .C0(n2368), .Y(n2370)
         );
  NAND3X2 U2198 ( .A(n2112), .B(n2111), .C(n2110), .Y(n2114) );
  NAND2XL U2199 ( .A(n2983), .B(\decoder/w_data_3[6] ), .Y(n2934) );
  NAND2XL U2200 ( .A(\decoder/w_data_3[7] ), .B(n2983), .Y(n2917) );
  NAND2XL U2201 ( .A(n2983), .B(\decoder/w_data_3[2] ), .Y(n2978) );
  NAND2XL U2202 ( .A(n2983), .B(\decoder/w_data_3[3] ), .Y(n2972) );
  NAND3X2 U2204 ( .A(n2905), .B(\decoder/w_PM_1[6] ), .C(\decoder/w_PM_2[6] ), 
        .Y(n2908) );
  OAI211X2 U2205 ( .A0(n2902), .A1(n2901), .B0(n2899), .C0(n2900), .Y(n1233)
         );
  NAND3X2 U2206 ( .A(n2853), .B(n2854), .C(n2852), .Y(n2857) );
  INVXL U2207 ( .A(n682), .Y(n2851) );
  NAND3X2 U2208 ( .A(n2861), .B(n2822), .C(n2862), .Y(n2831) );
  NAND2X2 U2209 ( .A(n2520), .B(n2521), .Y(n2514) );
  NAND2X2 U2210 ( .A(n2511), .B(n2531), .Y(n2509) );
  NAND2XL U2211 ( .A(n2489), .B(n2488), .Y(n2490) );
  NOR2X2 U2212 ( .A(n2485), .B(n2482), .Y(n2496) );
  XNOR2X4 U2213 ( .A(n2479), .B(n2478), .Y(n2520) );
  NAND2BX8 U2214 ( .AN(n344), .B(\decoder/w_enc_bit_8[0] ), .Y(n2432) );
  CLKAND2X4 U2216 ( .A(n2288), .B(n2293), .Y(n2294) );
  BUFX2 U2218 ( .A(n2391), .Y(n1614) );
  BUFX2 U2219 ( .A(n2394), .Y(n1619) );
  NOR2XL U2220 ( .A(n1786), .B(n1764), .Y(n929) );
  NAND3X2 U2222 ( .A(n2763), .B(n3095), .C(n2762), .Y(n2748) );
  NAND3X2 U2224 ( .A(n2759), .B(n1148), .C(n2758), .Y(n2762) );
  INVXL U2225 ( .A(n1148), .Y(n2791) );
  NAND3X2 U2228 ( .A(n2231), .B(n2232), .C(n2308), .Y(n2235) );
  NAND3X2 U2229 ( .A(n2232), .B(n2307), .C(n2229), .Y(n2236) );
  INVXL U2230 ( .A(n2647), .Y(n2649) );
  INVXL U2231 ( .A(n1734), .Y(n1747) );
  NOR2X2 U2232 ( .A(n2379), .B(n2375), .Y(n1281) );
  NAND3X2 U2233 ( .A(n1245), .B(n2192), .C(n2183), .Y(n2191) );
  NAND2X2 U2234 ( .A(n2177), .B(n2546), .Y(n2181) );
  INVXL U2235 ( .A(n2363), .Y(n2364) );
  OAI2BB1X2 U2236 ( .A0N(n2356), .A1N(n2357), .B0(n2360), .Y(n2348) );
  NAND2XL U2237 ( .A(n2260), .B(n2250), .Y(n2107) );
  NAND3X4 U2238 ( .A(n992), .B(n2915), .C(n2916), .Y(n2980) );
  INVXL U2239 ( .A(n668), .Y(n2898) );
  NAND3X2 U2240 ( .A(n2857), .B(n2856), .C(n2855), .Y(n2858) );
  NOR2XL U2241 ( .A(n1982), .B(n1980), .Y(n1942) );
  OAI2BB1X4 U2242 ( .A0N(n2283), .A1N(n2282), .B0(n2281), .Y(n2296) );
  NAND3X2 U2243 ( .A(n2280), .B(n2278), .C(n2279), .Y(n2281) );
  AOI2BB1X4 U2245 ( .A0N(n2636), .A1N(n2655), .B0(n1187), .Y(n2640) );
  NOR2BX2 U2246 ( .AN(\decoder/u_ACS_matrix/w_PM_6_to_7_1[2] ), .B(n2607), .Y(
        n1296) );
  INVXL U2247 ( .A(n1977), .Y(n1978) );
  NAND2XL U2248 ( .A(n1922), .B(n2937), .Y(n1923) );
  NAND3X2 U2249 ( .A(n1686), .B(n1774), .C(n1685), .Y(n1690) );
  INVXL U2250 ( .A(n2300), .Y(n2301) );
  NOR2XL U2251 ( .A(n1958), .B(n2939), .Y(n836) );
  NOR2XL U2252 ( .A(n2710), .B(n1097), .Y(n719) );
  INVXL U2253 ( .A(n2090), .Y(n2091) );
  INVXL U2256 ( .A(n1959), .Y(n1960) );
  INVXL U2257 ( .A(n2537), .Y(n2538) );
  OAI211X2 U2258 ( .A0(n2684), .A1(n2686), .B0(n2687), .C0(n2685), .Y(n1291)
         );
  NAND2XL U2259 ( .A(n2700), .B(n2699), .Y(n2689) );
  INVXL U2260 ( .A(n2315), .Y(n2316) );
  NAND3X2 U2261 ( .A(n2465), .B(n2464), .C(n2534), .Y(n2470) );
  NAND3X2 U2262 ( .A(n2465), .B(n2464), .C(n2460), .Y(n2462) );
  NAND3X2 U2263 ( .A(n2457), .B(n1605), .C(n2458), .Y(n2465) );
  NOR2XL U2267 ( .A(n1623), .B(n2968), .Y(n744) );
  NAND3X2 U2268 ( .A(n1285), .B(n1284), .C(n1281), .Y(n1267) );
  NAND3X2 U2269 ( .A(n2193), .B(n1282), .C(n1283), .Y(n1268) );
  NAND3X2 U2270 ( .A(n1283), .B(n1282), .C(n2380), .Y(n1266) );
  NAND3X2 U2271 ( .A(n2206), .B(n2191), .C(n2199), .Y(n1283) );
  NAND3X2 U2272 ( .A(n2208), .B(n1284), .C(n1285), .Y(n1265) );
  NAND3X2 U2273 ( .A(n2206), .B(n1261), .C(n2205), .Y(n1285) );
  NAND3BX2 U2274 ( .AN(n2178), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_4[0] ), 
        .C(n2177), .Y(n1244) );
  OAI2BB1X4 U2275 ( .A0N(n2037), .A1N(n2038), .B0(n2036), .Y(n2079) );
  OAI2BB1X4 U2276 ( .A0N(n1286), .A1N(n1815), .B0(n1816), .Y(n1820) );
  NAND2BX8 U2277 ( .AN(n328), .B(\decoder/w_enc_bit_4[0] ), .Y(n1893) );
  OAI2BB1X4 U2278 ( .A0N(n2374), .A1N(n2373), .B0(n2372), .Y(n2965) );
  NAND3X2 U2279 ( .A(n2878), .B(n2894), .C(n668), .Y(n2883) );
  NAND2XL U2280 ( .A(n2863), .B(n2881), .Y(n2802) );
  NAND2BX8 U2282 ( .AN(\decoder/w_enc_bit_6[0] ), .B(n1613), .Y(n2255) );
  NOR2XL U2283 ( .A(n2402), .B(n2401), .Y(n1116) );
  NOR2XL U2284 ( .A(n1187), .B(n2655), .Y(n733) );
  NOR2XL U2285 ( .A(n2784), .B(n2783), .Y(n666) );
  NOR2XL U2286 ( .A(n2953), .B(n1173), .Y(n846) );
  AOI21X2 U2287 ( .A0(n2718), .A1(n2717), .B0(n2772), .Y(n2769) );
  NAND2XL U2289 ( .A(n313), .B(\decoder/w_enc_bit_2[0] ), .Y(n1694) );
  OAI2BB1X2 U2290 ( .A0N(n2547), .A1N(n2565), .B0(n2548), .Y(n2575) );
  NAND3X2 U2291 ( .A(n2467), .B(n2468), .C(n2466), .Y(n2469) );
  NAND3X2 U2292 ( .A(n2467), .B(n2468), .C(n2452), .Y(n2463) );
  NAND3X2 U2293 ( .A(n2447), .B(n2454), .C(n2453), .Y(n2468) );
  NAND3X2 U2294 ( .A(n2441), .B(n2457), .C(n1605), .Y(n2467) );
  NAND3X2 U2295 ( .A(n2421), .B(n2422), .C(n2537), .Y(n2444) );
  NAND3X2 U2296 ( .A(n2197), .B(n2198), .C(n2381), .Y(n1282) );
  NAND3X2 U2297 ( .A(n2197), .B(n2198), .C(n1260), .Y(n1284) );
  NAND2XL U2298 ( .A(n994), .B(n2547), .Y(n2202) );
  NAND3X2 U2299 ( .A(n1776), .B(n1774), .C(n1775), .Y(n1226) );
  NAND3X2 U2300 ( .A(n1855), .B(n1854), .C(n1962), .Y(n1856) );
  INVXL U2301 ( .A(n1841), .Y(n1843) );
  INVXL U2302 ( .A(n2362), .Y(n2365) );
  NAND3X2 U2303 ( .A(n2348), .B(n2347), .C(n999), .Y(n2355) );
  NOR2XL U2304 ( .A(n2046), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_3[1] ), .Y(
        n2047) );
  OAI2BB1X2 U2305 ( .A0N(n1955), .A1N(n1933), .B0(n1945), .Y(n1951) );
  AOI21X2 U2306 ( .A0(n2285), .A1(n2284), .B0(n2324), .Y(n2312) );
  INVXL U2307 ( .A(n2264), .Y(n2266) );
  OAI2BB1X4 U2308 ( .A0N(n2640), .A1N(n2639), .B0(n2638), .Y(n2969) );
  BUFX2 U2309 ( .A(n3039), .Y(n1631) );
  BUFX2 U2310 ( .A(n3039), .Y(n1632) );
  BUFX2 U2311 ( .A(n3039), .Y(n1625) );
  BUFX2 U2312 ( .A(n3039), .Y(n1633) );
  BUFX2 U2314 ( .A(n3039), .Y(n1629) );
  BUFX2 U2315 ( .A(n3039), .Y(n1628) );
  BUFX2 U2316 ( .A(n3039), .Y(n1626) );
  BUFX2 U2317 ( .A(n3039), .Y(n1627) );
  BUFX2 U2318 ( .A(n3039), .Y(n1630) );
  NAND2XL U2319 ( .A(n1644), .B(n1645), .Y(n348) );
  CLKBUFX4 U2320 ( .A(n2392), .Y(n1617) );
  INVXL U2322 ( .A(n1708), .Y(n1760) );
  NOR2XL U2325 ( .A(n1127), .B(n2967), .Y(n731) );
  INVXL U2326 ( .A(n2551), .Y(n2554) );
  OAI2BB1X2 U2327 ( .A0N(n2544), .A1N(n2184), .B0(n2207), .Y(n2382) );
  OA21X2 U2328 ( .A0(\decoder/u_ACS_matrix/w_PM_3_to_4_4[1] ), .A1(n1866), 
        .B0(n1870), .Y(n1926) );
  NAND2X2 U2329 ( .A(n2086), .B(n1975), .Y(n2032) );
  NAND3X2 U2332 ( .A(n2473), .B(n2432), .C(
        \decoder/u_ACS_matrix/w_PM_7_to_8_2[0] ), .Y(n2471) );
  NAND2X2 U2333 ( .A(n1946), .B(n2088), .Y(n2051) );
  INVX2 U2334 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_3[6] ), .Y(n2798) );
  INVX2 U2335 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_3[4] ), .Y(n2930) );
  INVX2 U2336 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_3[3] ), .Y(n2946) );
  INVX2 U2337 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_3[2] ), .Y(n2957) );
  INVX2 U2338 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_3[5] ), .Y(n2793) );
  INVX2 U2339 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_3[5] ), .Y(n2933) );
  INVX2 U2340 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_3[4] ), .Y(n2949) );
  INVX2 U2341 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_3[3] ), .Y(n2961) );
  INVX2 U2342 ( .A(n1926), .Y(n1927) );
  INVX2 U2343 ( .A(n2303), .Y(n1328) );
  AND4X2 U2344 ( .A(n1649), .B(n1648), .C(n1647), .D(n1646), .Y(n311) );
  NAND2BX2 U2345 ( .AN(\decoder/u_input_shifter/U_input_split/N43 ), .B(n326), 
        .Y(n1496) );
  NAND2BX2 U2346 ( .AN(\decoder/u_input_shifter/U_input_split/N49 ), .B(n338), 
        .Y(n1355) );
  NAND2BX2 U2347 ( .AN(\decoder/u_input_shifter/U_input_split/N45 ), .B(n330), 
        .Y(n1540) );
  AND4X2 U2348 ( .A(n1653), .B(n1652), .C(n1651), .D(n1650), .Y(n318) );
  AND4X2 U2349 ( .A(n1657), .B(n1656), .C(n1655), .D(n1654), .Y(n315) );
  NOR2X2 U2350 ( .A(n1640), .B(n465), .Y(
        \decoder/u_input_shifter/u_input_fifo/N28 ) );
  AND4X2 U2351 ( .A(n1970), .B(n1969), .C(n1968), .D(n1967), .Y(n334) );
  NAND4X2 U2352 ( .A(n1974), .B(n1973), .C(n1972), .D(n1971), .Y(
        \decoder/u_input_shifter/U_input_split/N47 ) );
  NAND2BX2 U2353 ( .AN(n322), .B(\decoder/u_input_shifter/U_input_split/N41 ), 
        .Y(n1474) );
  NAND4X2 U2354 ( .A(n1675), .B(n1674), .C(n1673), .D(n1672), .Y(
        \decoder/u_input_shifter/U_input_split/N41 ) );
  AND4X2 U2355 ( .A(n1679), .B(n1678), .C(n1677), .D(n1676), .Y(n322) );
  NAND2BX2 U2356 ( .AN(n330), .B(\decoder/u_input_shifter/U_input_split/N45 ), 
        .Y(n1400) );
  NAND4X2 U2357 ( .A(n1832), .B(n1831), .C(n1830), .D(n1829), .Y(
        \decoder/u_input_shifter/U_input_split/N45 ) );
  AND4X2 U2358 ( .A(n1828), .B(n1827), .C(n1826), .D(n1825), .Y(n330) );
  NAND4X2 U2359 ( .A(n2399), .B(n2398), .C(n2397), .D(n2396), .Y(
        \decoder/u_input_shifter/U_input_split/N51 ) );
  NAND2BX2 U2360 ( .AN(n338), .B(\decoder/u_input_shifter/U_input_split/N49 ), 
        .Y(n1589) );
  NAND4X2 U2361 ( .A(n2140), .B(n2139), .C(n2138), .D(n2137), .Y(
        \decoder/u_input_shifter/U_input_split/N49 ) );
  AND4X2 U2362 ( .A(n2136), .B(n2135), .C(n2134), .D(n2133), .Y(n338) );
  NOR2X2 U2363 ( .A(n1645), .B(n1643), .Y(n2388) );
  NOR2X2 U2364 ( .A(n1644), .B(n347), .Y(n2395) );
  INVX2 U2365 ( .A(n1642), .Y(n1644) );
  INVX2 U2366 ( .A(n347), .Y(n1643) );
  INVX2 U2367 ( .A(n487), .Y(n2986) );
  NOR2X2 U2368 ( .A(n347), .B(n1645), .Y(n2394) );
  OR2X2 U2369 ( .A(n484), .B(n487), .Y(n1640) );
  NAND2X2 U2370 ( .A(n1670), .B(\decoder/u_ACS_matrix/w_PM_1_to_2_1[0] ), .Y(
        n1668) );
  NAND2X2 U2371 ( .A(n1670), .B(\decoder/u_ACS_matrix/w_PM_1_to_2_4[0] ), .Y(
        n1669) );
  INVX2 U2372 ( .A(n1667), .Y(n1670) );
  NAND2BX2 U2373 ( .AN(n465), .B(n487), .Y(n1636) );
  INVX2 U2374 ( .A(n465), .Y(n1639) );
  NAND2BX2 U2375 ( .AN(n1765), .B(n1773), .Y(n1685) );
  NAND2BX2 U2376 ( .AN(n1725), .B(n1724), .Y(n1686) );
  NAND2BX2 U2377 ( .AN(n1724), .B(n1725), .Y(n1688) );
  NAND2BX2 U2378 ( .AN(n1721), .B(n1722), .Y(n1689) );
  INVX2 U2379 ( .A(n1683), .Y(n1722) );
  NAND2X2 U2380 ( .A(n1684), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_3[1] ), .Y(
        n1683) );
  NAND2X2 U2381 ( .A(n1766), .B(n1772), .Y(n1684) );
  INVX2 U2382 ( .A(n1721), .Y(n1691) );
  INVX2 U2383 ( .A(n1687), .Y(n1721) );
  NAND2X2 U2384 ( .A(n1682), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_4[1] ), .Y(
        n1687) );
  NAND2X2 U2385 ( .A(n1767), .B(n1765), .Y(n1682) );
  INVX2 U2388 ( .A(\decoder/u_ACS_matrix/w_data_2_to_3_2[1] ), .Y(n1764) );
  NAND2BX2 U2390 ( .AN(n1728), .B(n1727), .Y(n1259) );
  NAND2X2 U2391 ( .A(n1726), .B(n1716), .Y(n1717) );
  INVX2 U2392 ( .A(n1720), .Y(n1726) );
  INVX2 U2393 ( .A(n1715), .Y(n1720) );
  NAND2X2 U2395 ( .A(n1710), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_1[1] ), .Y(
        n1719) );
  NAND2X2 U2396 ( .A(n1752), .B(n1760), .Y(n1710) );
  NOR2X2 U2397 ( .A(n1659), .B(n1658), .Y(n1661) );
  NAND2X2 U2398 ( .A(n1697), .B(n1694), .Y(n1660) );
  INVX2 U2399 ( .A(n1781), .Y(n1593) );
  NAND2X2 U2400 ( .A(n1729), .B(n1787), .Y(n1758) );
  INVX2 U2401 ( .A(n1784), .Y(n1757) );
  NAND2X2 U2402 ( .A(n1753), .B(n1760), .Y(n1756) );
  INVX2 U2403 ( .A(n1711), .Y(n1753) );
  NOR2X2 U2404 ( .A(n1713), .B(n1712), .Y(n1711) );
  INVX2 U2405 ( .A(\decoder/u_ACS_matrix/w_PM_2_to_3_2[0] ), .Y(n1712) );
  NAND2X2 U2406 ( .A(n1755), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_1[1] ), .Y(
        n1763) );
  NAND2X2 U2407 ( .A(n1752), .B(n1751), .Y(n1755) );
  XOR2X1 U2409 ( .A(n2749), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_4[5] ), .Y(
        n1174) );
  NAND2X2 U2411 ( .A(n2772), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[5] ), .Y(
        n2753) );
  NAND2X2 U2414 ( .A(n2718), .B(n2744), .Y(n2780) );
  NAND2X2 U2415 ( .A(n2714), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[3] ), .Y(
        n2718) );
  INVX2 U2416 ( .A(n2754), .Y(n2755) );
  INVX2 U2419 ( .A(n2741), .Y(n2788) );
  NAND2X2 U2420 ( .A(n2738), .B(n1299), .Y(n2740) );
  NAND2X2 U2423 ( .A(n2722), .B(n2737), .Y(n1301) );
  NAND2X2 U2426 ( .A(n2214), .B(n2302), .Y(n2216) );
  INVX2 U2428 ( .A(n2302), .Y(n2240) );
  NAND2X2 U2430 ( .A(n2328), .B(n2327), .Y(n2214) );
  INVX2 U2433 ( .A(n2217), .Y(n2212) );
  NAND2X2 U2435 ( .A(n2238), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_3[3] ), .Y(
        n2237) );
  INVX2 U2437 ( .A(n2230), .Y(n2231) );
  INVX2 U2439 ( .A(n2226), .Y(n2310) );
  NOR2X2 U2440 ( .A(n1163), .B(n1907), .Y(n1915) );
  OR2X2 U2441 ( .A(n1909), .B(n1908), .Y(n1163) );
  NOR2X2 U2442 ( .A(n1904), .B(n1905), .Y(n1907) );
  NAND2BX2 U2444 ( .AN(n3091), .B(n1897), .Y(n1899) );
  NOR2X2 U2447 ( .A(n2707), .B(n2706), .Y(n2682) );
  NAND2X2 U2448 ( .A(n2709), .B(n2664), .Y(n2680) );
  INVX2 U2449 ( .A(n2708), .Y(n2664) );
  INVX2 U2450 ( .A(n2670), .Y(n2709) );
  NAND2X2 U2453 ( .A(n2667), .B(n2787), .Y(n2739) );
  INVX2 U2457 ( .A(n2787), .Y(n2666) );
  INVX2 U2458 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_3[1] ), .Y(n2736) );
  INVX2 U2460 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_4[4] ), .Y(n1216) );
  INVX2 U2461 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_4[3] ), .Y(n1219) );
  NAND2X2 U2462 ( .A(n2676), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[3] ), .Y(
        n2673) );
  INVX2 U2463 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_3[6] ), .Y(n2752) );
  NAND3BX2 U2464 ( .AN(n2715), .B(n2676), .C(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[5] ), .Y(n2677) );
  NAND2X2 U2466 ( .A(n2722), .B(n2737), .Y(n1318) );
  NAND2X2 U2467 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_4[4] ), .B(
        \decoder/u_ACS_matrix/w_PM_7_to_8_4[3] ), .Y(n2659) );
  NAND2X2 U2468 ( .A(n1697), .B(n1696), .Y(n1698) );
  NAND2BX2 U2469 ( .AN(n1701), .B(n1700), .Y(n1693) );
  NAND2X2 U2470 ( .A(n1667), .B(\decoder/u_ACS_matrix/w_PM_1_to_2_3[0] ), .Y(
        n1695) );
  NAND2X2 U2471 ( .A(n1664), .B(n1666), .Y(n1667) );
  NAND2BX2 U2472 ( .AN(n2585), .B(n2584), .Y(n1280) );
  NAND2X2 U2473 ( .A(n2566), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[3] ), .Y(
        n2565) );
  NAND2BX2 U2475 ( .AN(n2548), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[5] ), 
        .Y(n2652) );
  NAND2BX2 U2476 ( .AN(n2551), .B(n1242), .Y(n2550) );
  NOR2X2 U2477 ( .A(n1316), .B(n1243), .Y(n1242) );
  INVX2 U2478 ( .A(n2533), .Y(n2466) );
  NOR2X2 U2480 ( .A(n2442), .B(n2436), .Y(n2440) );
  NAND2X2 U2482 ( .A(n2489), .B(n2484), .Y(n2433) );
  NAND2X2 U2483 ( .A(n2424), .B(n2435), .Y(n2425) );
  INVX2 U2485 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_1[5] ), .Y(n2450) );
  NAND2X2 U2486 ( .A(n2448), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_1[4] ), .Y(
        n2451) );
  INVX2 U2487 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_1[3] ), .Y(n2415) );
  NAND2BX2 U2490 ( .AN(n1838), .B(n1837), .Y(n1744) );
  INVX2 U2491 ( .A(n1742), .Y(n1837) );
  NAND2X2 U2492 ( .A(n1838), .B(n1742), .Y(n1741) );
  INVX2 U2494 ( .A(n1835), .Y(n1735) );
  NAND2BX2 U2495 ( .AN(n1734), .B(n1733), .Y(n1835) );
  NOR2X2 U2496 ( .A(n1736), .B(n1871), .Y(n1731) );
  NAND2X2 U2497 ( .A(n1737), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_4[1] ), .Y(
        n1736) );
  NAND2BX2 U2498 ( .AN(n1864), .B(n1862), .Y(n1737) );
  NOR2X2 U2499 ( .A(n1732), .B(n1865), .Y(n1734) );
  NAND2X2 U2500 ( .A(n1739), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_3[1] ), .Y(
        n1732) );
  INVX2 U2502 ( .A(\decoder/u_ACS_matrix/w_data_3_to_4_3[2] ), .Y(n1890) );
  INVX2 U2503 ( .A(\decoder/u_ACS_matrix/w_data_3_to_4_4[2] ), .Y(n1889) );
  NAND2X2 U2504 ( .A(n2194), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[5] ), .Y(
        n2375) );
  INVX2 U2505 ( .A(n2382), .Y(n2199) );
  NAND2X2 U2506 ( .A(n2192), .B(n1245), .Y(n2198) );
  NAND2X2 U2508 ( .A(n2192), .B(n2204), .Y(n1261) );
  INVX2 U2509 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_3[4] ), .Y(n2547) );
  NOR2X2 U2510 ( .A(n2380), .B(n2382), .Y(n2205) );
  NAND2BX2 U2512 ( .AN(n1602), .B(n1250), .Y(n2207) );
  OR2X2 U2513 ( .A(n2544), .B(n1601), .Y(n1602) );
  INVX2 U2514 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_4[4] ), .Y(n2544) );
  NAND2X2 U2515 ( .A(n2386), .B(n1251), .Y(n1270) );
  INVX2 U2516 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_3[1] ), .Y(n2171) );
  INVX2 U2518 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_4[3] ), .Y(n1601) );
  INVX2 U2519 ( .A(n1874), .Y(n1929) );
  INVX2 U2520 ( .A(n1930), .Y(n1883) );
  INVX2 U2521 ( .A(n1922), .Y(n1872) );
  NAND2X2 U2522 ( .A(n1867), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_3[1] ), .Y(
        n1868) );
  NAND2X2 U2523 ( .A(n1879), .B(n1880), .Y(n1888) );
  NOR2X2 U2525 ( .A(n1240), .B(\decoder/w_enc_bit_4[0] ), .Y(n1864) );
  INVX2 U2526 ( .A(n1875), .Y(n1879) );
  INVX2 U2527 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_4[2] ), .Y(n1871) );
  NAND2X2 U2528 ( .A(n1862), .B(n1882), .Y(n1866) );
  NAND2X2 U2530 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_4[0] ), .B(n1804), .Y(
        n1862) );
  INVX2 U2531 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_4[2] ), .Y(n2942) );
  INVX2 U2532 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_3[2] ), .Y(n2941) );
  NAND2X2 U2533 ( .A(n1778), .B(n1790), .Y(n1777) );
  INVX2 U2534 ( .A(n1771), .Y(n1790) );
  NAND2X2 U2535 ( .A(n1769), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_4[1] ), .Y(
        n1778) );
  NAND2BX2 U2536 ( .AN(n1797), .B(n1798), .Y(n1773) );
  NAND2BX2 U2537 ( .AN(n1798), .B(n1797), .Y(n1774) );
  NAND2X2 U2538 ( .A(n1767), .B(n1772), .Y(n1769) );
  OR2X2 U2539 ( .A(n324), .B(\decoder/w_enc_bit_3[0] ), .Y(n1772) );
  NAND2X2 U2540 ( .A(n1713), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_4[0] ), .Y(
        n1767) );
  NAND2X2 U2541 ( .A(n1766), .B(n1765), .Y(n1770) );
  NAND2X2 U2542 ( .A(n324), .B(\decoder/w_enc_bit_3[0] ), .Y(n1765) );
  NAND2X2 U2543 ( .A(n1713), .B(\decoder/u_ACS_matrix/w_PM_2_to_3_3[0] ), .Y(
        n1766) );
  OAI2B11X2 U2544 ( .A1N(n716), .A0(n2980), .B0(n2951), .C0(n2950), .Y(
        \decoder/u_cmp_sel/N47 ) );
  OAI2B11X2 U2545 ( .A1N(n717), .A0(n2980), .B0(n2963), .C0(n2962), .Y(
        \decoder/u_cmp_sel/N46 ) );
  INVX2 U2546 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_4[4] ), .Y(n2249) );
  INVX2 U2547 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_3[4] ), .Y(n2248) );
  INVX2 U2548 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_4[3] ), .Y(n2926) );
  INVX2 U2549 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_3[3] ), .Y(n2925) );
  INVX2 U2551 ( .A(n2082), .Y(n2028) );
  INVX2 U2552 ( .A(n2027), .Y(n2083) );
  NAND2X2 U2553 ( .A(n2076), .B(n2016), .Y(n2037) );
  NOR2X2 U2554 ( .A(n2021), .B(n2018), .Y(n1610) );
  INVX2 U2555 ( .A(n2077), .Y(n2016) );
  NAND2X2 U2556 ( .A(n2017), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_2[3] ), .Y(
        n2077) );
  NOR2X2 U2557 ( .A(n2021), .B(n2018), .Y(n2017) );
  NAND2BX2 U2559 ( .AN(n2013), .B(n1137), .Y(n2022) );
  INVX2 U2563 ( .A(\decoder/u_ACS_matrix/w_data_4_to_5_1[2] ), .Y(n2921) );
  INVX2 U2564 ( .A(\decoder/u_ACS_matrix/w_data_4_to_5_2[2] ), .Y(n2922) );
  INVX2 U2566 ( .A(n1957), .Y(n1596) );
  INVX2 U2567 ( .A(n1181), .Y(n1595) );
  INVX2 U2568 ( .A(n1963), .Y(n1854) );
  OR2X2 U2569 ( .A(n1849), .B(n2014), .Y(n1181) );
  NAND2X2 U2572 ( .A(n1841), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_2[1] ), .Y(
        n1851) );
  NAND2BX2 U2573 ( .AN(n2032), .B(n1846), .Y(n1847) );
  NAND2BX2 U2574 ( .AN(\decoder/u_ACS_matrix/w_PM_4_to_5_2[0] ), .B(
        \decoder/u_ACS_matrix/w_PM_4_to_5_1[0] ), .Y(n2030) );
  INVX2 U2575 ( .A(n2011), .Y(n2023) );
  INVX2 U2577 ( .A(\decoder/u_ACS_matrix/w_PM_4_to_5_1[1] ), .Y(n2010) );
  INVX2 U2579 ( .A(\decoder/u_ACS_matrix/w_PM_4_to_5_2[1] ), .Y(n1842) );
  NAND2BX2 U2580 ( .AN(n2013), .B(n1135), .Y(n1841) );
  NOR2X2 U2581 ( .A(n2993), .B(n1258), .Y(n2013) );
  INVX2 U2582 ( .A(\decoder/u_ACS_matrix/w_PM_4_to_5_2[0] ), .Y(n1258) );
  INVX2 U2583 ( .A(\decoder/u_ACS_matrix/w_data_4_to_5_1[3] ), .Y(n2040) );
  INVX2 U2584 ( .A(\decoder/u_ACS_matrix/w_data_4_to_5_2[3] ), .Y(n2041) );
  INVX2 U2585 ( .A(n1818), .Y(n1800) );
  NAND2BX2 U2586 ( .AN(\decoder/u_ACS_matrix/w_PM_3_to_4_1[2] ), .B(n1810), 
        .Y(n1811) );
  NAND2X2 U2588 ( .A(n1817), .B(n1818), .Y(n1286) );
  NAND2BX2 U2589 ( .AN(n1898), .B(n1231), .Y(n1801) );
  INVX2 U2590 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_1[0] ), .Y(n1799) );
  NOR2X2 U2591 ( .A(n1905), .B(n1612), .Y(n1185) );
  INVX2 U2592 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_1[1] ), .Y(n1612) );
  NAND2BX2 U2593 ( .AN(n1891), .B(n1897), .Y(n1802) );
  INVX2 U2594 ( .A(\decoder/u_ACS_matrix/w_data_3_to_4_2[2] ), .Y(n1913) );
  INVX2 U2595 ( .A(\decoder/u_ACS_matrix/w_data_3_to_4_1[2] ), .Y(n1912) );
  NAND4BX2 U2596 ( .AN(n2371), .B(n2369), .C(n2370), .D(n2374), .Y(n2372) );
  NAND2X2 U2597 ( .A(n2358), .B(n2405), .Y(n2368) );
  NOR2X2 U2598 ( .A(n2403), .B(n2350), .Y(n2371) );
  INVX2 U2599 ( .A(n2404), .Y(n2350) );
  NAND2BX2 U2602 ( .AN(n2409), .B(n2339), .Y(n2357) );
  NAND2X2 U2603 ( .A(n2339), .B(n2410), .Y(n2356) );
  NAND2BX2 U2604 ( .AN(\decoder/u_ACS_matrix/w_PM_6_to_7_1[2] ), .B(n2335), 
        .Y(n2336) );
  NAND2X2 U2607 ( .A(n2330), .B(n2402), .Y(n2374) );
  INVX2 U2608 ( .A(n2353), .Y(n2402) );
  NAND2X2 U2609 ( .A(n2599), .B(n1155), .Y(n2331) );
  INVX2 U2610 ( .A(n2401), .Y(n2330) );
  NOR2X2 U2611 ( .A(n1095), .B(n1197), .Y(n1193) );
  INVX2 U2612 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_2[4] ), .Y(n1197) );
  INVX2 U2617 ( .A(n2125), .Y(n2156) );
  NAND2X2 U2618 ( .A(n2122), .B(n2121), .Y(n2125) );
  INVX2 U2621 ( .A(n2121), .Y(n2118) );
  NAND2BX2 U2622 ( .AN(n2132), .B(n2131), .Y(n2110) );
  INVX2 U2623 ( .A(n2109), .Y(n2131) );
  NAND2X2 U2624 ( .A(n2132), .B(n2109), .Y(n2108) );
  NAND2X2 U2627 ( .A(n2257), .B(n3025), .Y(n2116) );
  NAND2BX2 U2629 ( .AN(n1274), .B(n1273), .Y(n1986) );
  INVX2 U2630 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_4[1] ), .Y(n2220) );
  NOR2X2 U2631 ( .A(n2144), .B(n2143), .Y(n1995) );
  NOR2X2 U2632 ( .A(n2218), .B(n1606), .Y(n1183) );
  INVX2 U2633 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_3[3] ), .Y(n1606) );
  OAI2B11X2 U2634 ( .A1N(n715), .A0(n2980), .B0(n2935), .C0(n2934), .Y(
        \decoder/u_cmp_sel/N48 ) );
  OAI2B11X2 U2635 ( .A1N(n714), .A0(n2980), .B0(n2918), .C0(n2917), .Y(
        \decoder/u_cmp_sel/N49 ) );
  OAI2B11X2 U2636 ( .A1N(\decoder/w_data_1[2] ), .A0(n2980), .B0(n2979), .C0(
        n2978), .Y(\decoder/u_cmp_sel/N44 ) );
  OAI2B11X2 U2637 ( .A1N(n718), .A0(n2980), .B0(n2973), .C0(n2972), .Y(
        \decoder/u_cmp_sel/N45 ) );
  AOI2BB2X2 U2639 ( .B0(n2885), .B1(\decoder/w_PM_4[6] ), .A0N(n2884), .A1N(
        n682), .Y(n2911) );
  NAND2X2 U2640 ( .A(n2882), .B(n2881), .Y(n2907) );
  OR2X2 U2642 ( .A(n2873), .B(n2880), .Y(n2874) );
  OAI2B11X2 U2643 ( .A1N(n2891), .A0(n2870), .B0(n2868), .C0(n2867), .Y(n2875)
         );
  NAND2BX2 U2645 ( .AN(n2863), .B(n668), .Y(n2884) );
  INVX2 U2646 ( .A(\decoder/w_PM_2[6] ), .Y(n2872) );
  INVX2 U2647 ( .A(n2840), .Y(n2843) );
  INVX2 U2648 ( .A(n2836), .Y(n2833) );
  NAND2BX2 U2649 ( .AN(\decoder/w_PM_2[5] ), .B(\decoder/w_PM_1[5] ), .Y(n2836) );
  INVX2 U2650 ( .A(\decoder/w_PM_1[6] ), .Y(n2895) );
  NOR2X2 U2651 ( .A(n668), .B(n2845), .Y(n2866) );
  INVX2 U2652 ( .A(n695), .Y(n2845) );
  NAND2BX2 U2653 ( .AN(n2826), .B(n2825), .Y(n2852) );
  INVX2 U2654 ( .A(n697), .Y(n2834) );
  INVX2 U2655 ( .A(n699), .Y(n2864) );
  NAND2BX2 U2656 ( .AN(n1559), .B(n2821), .Y(n2861) );
  NAND2BX2 U2657 ( .AN(n685), .B(\decoder/w_PM_1[1] ), .Y(n2811) );
  NAND3BX2 U2658 ( .AN(n2807), .B(n2806), .C(n2809), .Y(n2814) );
  NAND2BX2 U2659 ( .AN(\decoder/w_PM_1[3] ), .B(n683), .Y(n2809) );
  INVX2 U2660 ( .A(n711), .Y(n2892) );
  NAND2BX2 U2661 ( .AN(\decoder/w_PM_1[5] ), .B(n681), .Y(n2808) );
  NAND2BX2 U2662 ( .AN(\decoder/w_PM_3[6] ), .B(\decoder/w_PM_1[6] ), .Y(n2804) );
  NAND2BX2 U2663 ( .AN(n681), .B(\decoder/w_PM_1[5] ), .Y(n2805) );
  NAND4BX2 U2664 ( .AN(n695), .B(n2828), .C(n682), .D(n2827), .Y(n2856) );
  NAND2BX2 U2665 ( .AN(\decoder/w_PM_2[6] ), .B(\decoder/w_PM_3[6] ), .Y(n2855) );
  NAND2BX2 U2666 ( .AN(\decoder/w_PM_3[6] ), .B(\decoder/w_PM_2[6] ), .Y(n2827) );
  NAND2BX2 U2667 ( .AN(\decoder/w_PM_3[6] ), .B(\decoder/w_PM_4[6] ), .Y(n2881) );
  INVX2 U2668 ( .A(\decoder/w_PM_3[6] ), .Y(n2906) );
  NAND2X2 U2669 ( .A(n1383), .B(n1381), .Y(n2976) );
  INVX2 U2670 ( .A(n2099), .Y(n2062) );
  NAND2X2 U2673 ( .A(n2053), .B(n2093), .Y(n2054) );
  INVX2 U2674 ( .A(n2052), .Y(n2093) );
  NAND2BX2 U2675 ( .AN(n2051), .B(n2067), .Y(n2055) );
  NAND2X2 U2676 ( .A(n2094), .B(n2052), .Y(n2067) );
  INVX2 U2678 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_1[5] ), .Y(n2929) );
  INVX2 U2679 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_1[3] ), .Y(n2956) );
  INVX2 U2680 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_1[6] ), .Y(n2792) );
  INVX2 U2681 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_1[2] ), .Y(n2966) );
  OR2X2 U2682 ( .A(n2974), .B(n1546), .Y(n1182) );
  INVX2 U2683 ( .A(n2511), .Y(n2532) );
  NAND2BX2 U2684 ( .AN(n2517), .B(n2516), .Y(n2508) );
  INVX2 U2685 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_2[5] ), .Y(n2505) );
  NAND2X2 U2686 ( .A(n2477), .B(n2472), .Y(n2517) );
  NAND2X2 U2687 ( .A(n1307), .B(n1207), .Y(n2472) );
  INVX2 U2688 ( .A(n1310), .Y(n1597) );
  NAND2X2 U2689 ( .A(n2498), .B(n2540), .Y(n2499) );
  INVX2 U2690 ( .A(n2497), .Y(n2540) );
  NAND2BX2 U2691 ( .AN(n1306), .B(n2481), .Y(n1307) );
  NAND2BX2 U2692 ( .AN(n2526), .B(n1139), .Y(n2493) );
  NOR2X2 U2694 ( .A(n2484), .B(n956), .Y(n2487) );
  INVX2 U2695 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_2[6] ), .Y(n2478) );
  NAND2X2 U2696 ( .A(n2506), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_2[5] ), .Y(
        n2479) );
  NOR2X2 U2698 ( .A(n1306), .B(n1207), .Y(n1208) );
  INVX2 U2699 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_2[4] ), .Y(n1207) );
  NAND2X2 U2700 ( .A(n748), .B(n749), .Y(n1306) );
  NAND2X2 U2701 ( .A(n2471), .B(n1204), .Y(n1220) );
  NAND2X2 U2702 ( .A(n2507), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_1[5] ), .Y(
        n2476) );
  INVX2 U2703 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_1[4] ), .Y(n2945) );
  INVX2 U2704 ( .A(\decoder/u_ACS_matrix/w_data_4_to_5_3[2] ), .Y(n2923) );
  INVX2 U2705 ( .A(\decoder/u_ACS_matrix/w_data_4_to_5_4[2] ), .Y(n2924) );
  NAND2X2 U2706 ( .A(n1138), .B(n1977), .Y(n1953) );
  NAND2X2 U2707 ( .A(n1951), .B(n1950), .Y(n1954) );
  INVX2 U2708 ( .A(n1946), .Y(n2089) );
  NAND2X2 U2709 ( .A(n967), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_3[3] ), .Y(
        n1952) );
  NAND2X2 U2710 ( .A(n1937), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_4[2] ), .Y(
        n1936) );
  INVX2 U2711 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_2[3] ), .Y(n2927) );
  INVX2 U2712 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_1[3] ), .Y(n2928) );
  INVX2 U2713 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_2[4] ), .Y(n2298) );
  INVX2 U2714 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_1[4] ), .Y(n2299) );
  INVX2 U2715 ( .A(n2288), .Y(n2325) );
  INVX2 U2716 ( .A(n2294), .Y(n2295) );
  NOR2X2 U2717 ( .A(n2294), .B(n2291), .Y(n2292) );
  INVX2 U2719 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_2[3] ), .Y(n2286) );
  INVX2 U2720 ( .A(n2293), .Y(n2324) );
  NAND2X2 U2721 ( .A(n1290), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[4] ), .Y(
        n2293) );
  INVX2 U2723 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_1[4] ), .Y(n2285) );
  AOI2BB2X2 U2725 ( .B0(n2271), .B1(n2270), .A0N(n2266), .A1N(n2265), .Y(n2274) );
  NAND2BX2 U2726 ( .AN(\decoder/u_ACS_matrix/w_PM_5_to_6_2[0] ), .B(
        \decoder/u_ACS_matrix/w_PM_5_to_6_1[0] ), .Y(n2260) );
  NAND2X2 U2727 ( .A(n1136), .B(n2321), .Y(n2263) );
  NAND2X2 U2728 ( .A(n2251), .B(n2254), .Y(n2264) );
  INVX2 U2729 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_2[1] ), .Y(n2256) );
  INVX2 U2730 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_2[2] ), .Y(n2943) );
  INVX2 U2731 ( .A(\decoder/u_ACS_matrix/w_data_5_to_6_1[2] ), .Y(n2944) );
  INVX2 U2732 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_1[3] ), .Y(n2948) );
  INVX2 U2733 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_1[5] ), .Y(n2795) );
  INVX2 U2734 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_1[4] ), .Y(n2932) );
  NAND2X2 U2736 ( .A(n2619), .B(n2618), .Y(n2643) );
  INVX2 U2737 ( .A(n2614), .Y(n2615) );
  INVX2 U2740 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_1[2] ), .Y(n2602) );
  INVX2 U2741 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_1[4] ), .Y(n2590) );
  OR2X2 U2742 ( .A(n1229), .B(n2594), .Y(n1187) );
  INVX2 U2745 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_1[5] ), .Y(n2593) );
  NAND2X2 U2746 ( .A(n2591), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_1[4] ), .Y(
        n1297) );
  INVX2 U2747 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_1[3] ), .Y(n2607) );
  INVX2 U2748 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_1[1] ), .Y(n2598) );
  NAND2X2 U2749 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_1[0] ), .B(n2604), .Y(
        n2589) );
  INVX2 U2750 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_1[2] ), .Y(n2959) );
  INVX2 U2751 ( .A(\decoder/u_ACS_matrix/w_data_6_to_7_2[2] ), .Y(n2960) );
  XNOR2X1 U2752 ( .A(n317), .B(n320), .Y(n2985) );
  NOR3X1 U2753 ( .A(n350), .B(n2986), .C(n1643), .Y(n2392) );
  NOR3BX1 U2754 ( .AN(n350), .B(n347), .C(n487), .Y(n2391) );
  NOR3X1 U2755 ( .A(n350), .B(n347), .C(n2986), .Y(n2390) );
  NAND2X2 U2756 ( .A(n350), .B(n487), .Y(n1645) );
  AND2X2 U2757 ( .A(n1642), .B(n347), .Y(n2389) );
  NOR2X2 U2758 ( .A(n350), .B(n487), .Y(n1642) );
  OAI21X1 U2759 ( .A0(n1670), .A1(\decoder/u_ACS_matrix/w_PM_1_to_2_4[0] ), 
        .B0(n1669), .Y(n1703) );
  XNOR2X1 U2760 ( .A(n2772), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[5] ), .Y(
        n2785) );
  OAI21X1 U2761 ( .A0(n2238), .A1(\decoder/u_ACS_matrix/w_PM_5_to_6_3[3] ), 
        .B0(n2237), .Y(n2304) );
  OAI21X1 U2762 ( .A0(n1667), .A1(\decoder/u_ACS_matrix/w_PM_1_to_2_3[0] ), 
        .B0(n1695), .Y(n1700) );
  NAND2BX2 U2763 ( .AN(\decoder/w_enc_bit_2[0] ), .B(n313), .Y(n1666) );
  NAND2BX2 U2764 ( .AN(n313), .B(\decoder/w_enc_bit_2[0] ), .Y(n1664) );
  INVX2 U2765 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_3[2] ), .Y(n2549) );
  OAI21X1 U2767 ( .A0(\decoder/u_ACS_matrix/w_PM_3_to_4_3[1] ), .A1(n1867), 
        .B0(n1868), .Y(n1928) );
  INVX2 U2768 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_3[2] ), .Y(n1865) );
  BUFX2 U2769 ( .A(n328), .Y(n1240) );
  INVX2 U2770 ( .A(\decoder/u_ACS_matrix/w_PM_4_to_5_2[2] ), .Y(n2018) );
  INVX2 U2771 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_1[2] ), .Y(n1905) );
  INVX2 U2773 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_3[2] ), .Y(n2218) );
  NAND2X2 U2774 ( .A(n1550), .B(n1548), .Y(n2974) );
  XNOR2X1 U2775 ( .A(n2993), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_3[0] ), .Y(
        n2088) );
  INVX2 U2776 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_1[2] ), .Y(n2270) );
  NOR2BX1 U2777 ( .AN(n2376), .B(n2375), .Y(n745) );
  NOR2BX1 U2778 ( .AN(n1072), .B(n2652), .Y(n720) );
  AOI22XL U2779 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_7[3] ), .B0(
        n1619), .B1(\decoder/u_input_shifter/w_data_4[3] ), .Y(n1646) );
  AOI22XL U2780 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_1[3] ), .B0(
        n1617), .B1(\decoder/u_input_shifter/w_data_2[3] ), .Y(n1647) );
  AOI22XL U2781 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_3[3] ), .B0(
        n1616), .B1(\decoder/u_input_shifter/w_data_8[3] ), .Y(n1648) );
  AOI22XL U2782 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_5[3] ), .B0(
        n1615), .B1(\decoder/u_input_shifter/w_data_6[3] ), .Y(n1649) );
  AOI22XL U2783 ( .A0(n1619), .A1(\decoder/u_input_shifter/w_data_5[1] ), .B0(
        n1616), .B1(\decoder/u_input_shifter/w_data_1[1] ), .Y(n1650) );
  AOI22XL U2784 ( .A0(n1615), .A1(\decoder/u_input_shifter/w_data_7[1] ), .B0(
        n1617), .B1(\decoder/u_input_shifter/w_data_3[1] ), .Y(n1651) );
  AOI22XL U2785 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_2[1] ), .B0(
        n1614), .B1(\decoder/u_input_shifter/w_data_6[1] ), .Y(n1652) );
  AOI22XL U2786 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_4[1] ), .B0(
        n1618), .B1(\decoder/u_input_shifter/w_data_8[1] ), .Y(n1653) );
  AOI22XL U2787 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_8[0] ), .B0(
        n1616), .B1(\decoder/u_input_shifter/w_data_1[0] ), .Y(n1654) );
  AOI22XL U2788 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_6[0] ), .B0(
        n1617), .B1(\decoder/u_input_shifter/w_data_3[0] ), .Y(n1655) );
  AOI22XL U2789 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_2[0] ), .B0(
        n1615), .B1(\decoder/u_input_shifter/w_data_7[0] ), .Y(n1656) );
  AOI22XL U2790 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_4[0] ), .B0(
        n1619), .B1(\decoder/u_input_shifter/w_data_5[0] ), .Y(n1657) );
  XNOR2X1 U2791 ( .A(\decoder/u_input_shifter/U_input_split/N47 ), .B(n334), 
        .Y(n1587) );
  AOI22XL U2792 ( .A0(n1619), .A1(\decoder/u_input_shifter/w_data_8[11] ), 
        .B0(n1616), .B1(\decoder/u_input_shifter/w_data_4[11] ), .Y(n1967) );
  AOI22XL U2793 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_1[11] ), 
        .B0(n1617), .B1(\decoder/u_input_shifter/w_data_6[11] ), .Y(n1968) );
  AOI22XL U2794 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_5[11] ), 
        .B0(n1615), .B1(\decoder/u_input_shifter/w_data_2[11] ), .Y(n1969) );
  AOI22XL U2795 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_7[11] ), 
        .B0(n1618), .B1(\decoder/u_input_shifter/w_data_3[11] ), .Y(n1970) );
  AOI22XL U2796 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_3[10] ), 
        .B0(n1619), .B1(\decoder/u_input_shifter/w_data_8[10] ), .Y(n1971) );
  AOI22XL U2797 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_5[10] ), 
        .B0(n1617), .B1(\decoder/u_input_shifter/w_data_6[10] ), .Y(n1972) );
  AOI22XL U2798 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_1[10] ), 
        .B0(n1615), .B1(\decoder/u_input_shifter/w_data_2[10] ), .Y(n1973) );
  AOI22XL U2799 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_7[10] ), 
        .B0(n1616), .B1(\decoder/u_input_shifter/w_data_4[10] ), .Y(n1974) );
  AOI22XL U2800 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_6[4] ), .B0(
        n1619), .B1(\decoder/u_input_shifter/w_data_3[4] ), .Y(n1672) );
  AOI22XL U2801 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_8[4] ), .B0(
        n1617), .B1(\decoder/u_input_shifter/w_data_1[4] ), .Y(n1673) );
  AOI22XL U2802 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_4[4] ), .B0(
        n1615), .B1(\decoder/u_input_shifter/w_data_5[4] ), .Y(n1674) );
  AOI22XL U2803 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_2[4] ), .B0(
        n1616), .B1(\decoder/u_input_shifter/w_data_7[4] ), .Y(n1675) );
  AOI22XL U2804 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_6[5] ), .B0(
        n1619), .B1(\decoder/u_input_shifter/w_data_3[5] ), .Y(n1676) );
  AOI22XL U2805 ( .A0(n1615), .A1(\decoder/u_input_shifter/w_data_5[5] ), .B0(
        n1617), .B1(\decoder/u_input_shifter/w_data_1[5] ), .Y(n1677) );
  AOI22XL U2806 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_8[5] ), .B0(
        n1614), .B1(\decoder/u_input_shifter/w_data_4[5] ), .Y(n1678) );
  AOI22XL U2807 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_2[5] ), .B0(
        n1616), .B1(\decoder/u_input_shifter/w_data_7[5] ), .Y(n1679) );
  AOI21X1 U2808 ( .A0(n1723), .A1(n1691), .B0(n1683), .Y(n900) );
  AOI22XL U2809 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_4[8] ), .B0(
        n1619), .B1(\decoder/u_input_shifter/w_data_1[8] ), .Y(n1829) );
  AOI22XL U2810 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_6[8] ), .B0(
        n1617), .B1(\decoder/u_input_shifter/w_data_7[8] ), .Y(n1830) );
  AOI22XL U2811 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_2[8] ), .B0(
        n1615), .B1(\decoder/u_input_shifter/w_data_3[8] ), .Y(n1831) );
  AOI22XL U2812 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_8[8] ), .B0(
        n1616), .B1(\decoder/u_input_shifter/w_data_5[8] ), .Y(n1832) );
  AOI22XL U2813 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_4[9] ), .B0(
        n1619), .B1(\decoder/u_input_shifter/w_data_1[9] ), .Y(n1825) );
  AOI22XL U2814 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_2[9] ), .B0(
        n1617), .B1(\decoder/u_input_shifter/w_data_7[9] ), .Y(n1826) );
  AOI22XL U2815 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_6[9] ), .B0(
        n1615), .B1(\decoder/u_input_shifter/w_data_3[9] ), .Y(n1827) );
  AOI22XL U2816 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_8[9] ), .B0(
        n1616), .B1(\decoder/u_input_shifter/w_data_5[9] ), .Y(n1828) );
  XNOR2X1 U2817 ( .A(\decoder/u_input_shifter/U_input_split/N51 ), .B(n342), 
        .Y(n1571) );
  AOI22XL U2818 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_1[14] ), 
        .B0(n1619), .B1(\decoder/u_input_shifter/w_data_6[14] ), .Y(n2396) );
  AOI22XL U2819 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_3[14] ), 
        .B0(n1617), .B1(\decoder/u_input_shifter/w_data_4[14] ), .Y(n2397) );
  AOI22XL U2820 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_7[14] ), 
        .B0(n1615), .B1(\decoder/u_input_shifter/w_data_8[14] ), .Y(n2398) );
  AOI22XL U2821 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_5[14] ), 
        .B0(n1616), .B1(\decoder/u_input_shifter/w_data_2[14] ), .Y(n2399) );
  AOI22XL U2822 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_2[12] ), 
        .B0(n1619), .B1(\decoder/u_input_shifter/w_data_7[12] ), .Y(n2137) );
  AOI22XL U2823 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_4[12] ), 
        .B0(n1617), .B1(\decoder/u_input_shifter/w_data_5[12] ), .Y(n2138) );
  AOI22XL U2824 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_8[12] ), 
        .B0(n1615), .B1(\decoder/u_input_shifter/w_data_1[12] ), .Y(n2139) );
  AOI22XL U2825 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_6[12] ), 
        .B0(n1616), .B1(\decoder/u_input_shifter/w_data_3[12] ), .Y(n2140) );
  AOI22XL U2826 ( .A0(n1618), .A1(\decoder/u_input_shifter/w_data_2[13] ), 
        .B0(n1616), .B1(\decoder/u_input_shifter/w_data_3[13] ), .Y(n2133) );
  AOI22XL U2827 ( .A0(n1614), .A1(\decoder/u_input_shifter/w_data_8[13] ), 
        .B0(n1617), .B1(\decoder/u_input_shifter/w_data_5[13] ), .Y(n2134) );
  AOI22XL U2828 ( .A0(n2393), .A1(\decoder/u_input_shifter/w_data_4[13] ), 
        .B0(n1615), .B1(\decoder/u_input_shifter/w_data_1[13] ), .Y(n2135) );
  AND3X2 U2829 ( .A(n2986), .B(n347), .C(n350), .Y(n2393) );
  AOI22XL U2830 ( .A0(n2389), .A1(\decoder/u_input_shifter/w_data_6[13] ), 
        .B0(n1619), .B1(\decoder/u_input_shifter/w_data_7[13] ), .Y(n2136) );
  NOR3BX1 U2831 ( .AN(n484), .B(n465), .C(n487), .Y(n951) );
  NAND2XL U2832 ( .A(n465), .B(n487), .Y(n1638) );
  MXI2X1 U2833 ( .A(n1703), .B(n1702), .S0(n1671), .Y(n936) );
  MXI2X1 U2834 ( .A(n1665), .B(n1164), .S0(n1671), .Y(n935) );
  AND2X2 U2835 ( .A(n1668), .B(n1666), .Y(n1164) );
  AND2X2 U2837 ( .A(n1669), .B(n1666), .Y(n1188) );
  MXI2X1 U2838 ( .A(n1700), .B(n1701), .S0(n1681), .Y(n932) );
  NOR3X1 U2839 ( .A(n487), .B(n1637), .C(n1639), .Y(n953) );
  MXI2X1 U2840 ( .A(n1798), .B(n971), .S0(n2919), .Y(n902) );
  MXI2X1 U2842 ( .A(n1701), .B(n1700), .S0(n1699), .Y(n939) );
  OAI2BB1X1 U2843 ( .A0N(n1731), .A1N(n1834), .B0(n1833), .Y(n880) );
  NAND2XL U2844 ( .A(n2936), .B(n1734), .Y(n1833) );
  MXI2X1 U2847 ( .A(n1929), .B(n1930), .S0(n2936), .Y(n883) );
  MXI2X1 U2849 ( .A(n1838), .B(n1837), .S0(n2936), .Y(n882) );
  OAI2BB1X1 U2850 ( .A0N(n1925), .A1N(n1924), .B0(n1923), .Y(n862) );
  OAI21X1 U2851 ( .A0(n1684), .A1(\decoder/u_ACS_matrix/w_PM_2_to_3_3[1] ), 
        .B0(n1683), .Y(n1724) );
  MXI2X1 U2852 ( .A(n1836), .B(n1835), .S0(n2936), .Y(n881) );
  AOI21X1 U2854 ( .A0(n1958), .A1(n1181), .B0(n1596), .Y(n829) );
  AOI21X1 U2855 ( .A0(n1793), .A1(n1771), .B0(n1792), .Y(n917) );
  MXI2X1 U2856 ( .A(n2701), .B(n2700), .S0(n1624), .Y(n694) );
  MXI2X1 U2857 ( .A(n2302), .B(n2301), .S0(n2964), .Y(n1114) );
  AND2X2 U2858 ( .A(n1720), .B(n1719), .Y(n1192) );
  OAI21X1 U2859 ( .A0(n1710), .A1(\decoder/u_ACS_matrix/w_PM_2_to_3_1[1] ), 
        .B0(n1719), .Y(n1728) );
  OAI21X1 U2860 ( .A0(n1693), .A1(n1680), .B0(n1594), .Y(n1663) );
  MXI2X1 U2864 ( .A(n2650), .B(n2651), .S0(n1120), .Y(n764) );
  OAI21X1 U2870 ( .A0(n2940), .A1(n2081), .B0(n2080), .Y(n851) );
  OAI21X1 U2872 ( .A0(n1755), .A1(\decoder/u_ACS_matrix/w_PM_2_to_3_1[1] ), 
        .B0(n1763), .Y(n1784) );
  AND3X2 U2878 ( .A(n2745), .B(n2779), .C(n2781), .Y(n2754) );
  MXI2X1 U2879 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_3[1] ), .B(n2736), .S0(
        n2735), .Y(n2789) );
  MXI2X1 U2882 ( .A(n2310), .B(n2311), .S0(n1620), .Y(n776) );
  OAI21X1 U2883 ( .A0(n2242), .A1(\decoder/u_ACS_matrix/w_PM_5_to_6_4[4] ), 
        .B0(n2215), .Y(n2302) );
  XNOR2X1 U2889 ( .A(n1909), .B(n1908), .Y(n1917) );
  AND2X2 U2890 ( .A(n1907), .B(n1163), .Y(n1190) );
  BUFX2 U2892 ( .A(n1893), .Y(n1231) );
  XNOR2X1 U2906 ( .A(n2673), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[4] ), .Y(
        n2690) );
  MXI2X1 U2910 ( .A(n974), .B(n2581), .S0(n1127), .Y(n723) );
  AND2X2 U2914 ( .A(n1695), .B(n1694), .Y(n1186) );
  NOR2BX1 U2915 ( .AN(n1701), .B(n1700), .Y(n1692) );
  XNOR2X1 U2917 ( .A(n1598), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[5] ), .Y(
        n2653) );
  OAI21X1 U2919 ( .A0(n2566), .A1(\decoder/u_ACS_matrix/w_PM_6_to_7_3[3] ), 
        .B0(n2565), .Y(n2581) );
  OAI21X1 U2920 ( .A0(\decoder/u_ACS_matrix/w_PM_6_to_7_4[3] ), .A1(n2564), 
        .B0(n2563), .Y(n2582) );
  OAI21X1 U2921 ( .A0(n2552), .A1(\decoder/u_ACS_matrix/w_PM_6_to_7_4[2] ), 
        .B0(n2550), .Y(n2585) );
  AOI21X1 U2922 ( .A0(n2549), .A1(n2555), .B0(n2566), .Y(n2583) );
  AND2X2 U2924 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_3[4] ), .B(
        \decoder/u_ACS_matrix/w_PM_6_to_7_3[3] ), .Y(n1315) );
  OAI21X1 U2927 ( .A0(\decoder/u_ACS_matrix/w_PM_7_to_8_2[1] ), .A1(n2431), 
        .B0(n2430), .Y(n2530) );
  MXI2X1 U2933 ( .A(n1889), .B(n1890), .S0(n2936), .Y(n884) );
  XNOR2X1 U2934 ( .A(n1739), .B(n1738), .Y(n1742) );
  OAI21X1 U2935 ( .A0(n1737), .A1(\decoder/u_ACS_matrix/w_PM_3_to_4_4[1] ), 
        .B0(n1736), .Y(n1838) );
  XNOR2X1 U2937 ( .A(n1736), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_4[2] ), .Y(
        n1743) );
  NOR2BX1 U2939 ( .AN(n2202), .B(n2201), .Y(n2183) );
  NAND2XL U2940 ( .A(n2983), .B(n1462), .Y(n2984) );
  AOI21X1 U2941 ( .A0(n1883), .A1(n1929), .B0(n1882), .Y(n1884) );
  OAI21X1 U2942 ( .A0(n1881), .A1(n1878), .B0(n1877), .Y(n1887) );
  OAI21X1 U2944 ( .A0(n1713), .A1(\decoder/u_ACS_matrix/w_PM_2_to_3_4[0] ), 
        .B0(n1767), .Y(n1798) );
  XNOR2X1 U2945 ( .A(n1769), .B(n1768), .Y(n1794) );
  OAI21X1 U2949 ( .A0(\decoder/u_ACS_matrix/w_PM_4_to_5_2[1] ), .A1(n2022), 
        .B0(n2021), .Y(n2085) );
  AOI21X1 U2950 ( .A0(n2018), .A1(n2021), .B0(n1610), .Y(n2027) );
  XNOR2X1 U2954 ( .A(n1851), .B(n2018), .Y(n1963) );
  XNOR2X1 U2956 ( .A(\decoder/u_ACS_matrix/w_PM_4_to_5_2[0] ), .B(n2993), .Y(
        n1975) );
  OAI21X1 U2957 ( .A0(\decoder/u_ACS_matrix/w_PM_4_to_5_1[0] ), .A1(n1845), 
        .B0(n2025), .Y(n2086) );
  OAI2BB1X1 U2960 ( .A0N(n1806), .A1N(n1895), .B0(n1896), .Y(n1808) );
  AOI21X1 U2967 ( .A0(n2401), .A1(n2353), .B0(n2352), .Y(n2354) );
  AND2X2 U2969 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_1[1] ), .B(
        \decoder/u_ACS_matrix/w_PM_6_to_7_1[2] ), .Y(n1239) );
  OAI2BB1X1 U2973 ( .A0N(n2106), .A1N(n2252), .B0(n2105), .Y(n2132) );
  XNOR2X1 U2974 ( .A(n2116), .B(n2256), .Y(n2109) );
  AND3X2 U2977 ( .A(n1997), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_4[1] ), .C(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[3] ), .Y(n1273) );
  XNOR2X1 U2980 ( .A(n2211), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_3[0] ), .Y(
        n2226) );
  OAI21X1 U2983 ( .A0(n2905), .A1(\decoder/w_PM_2[6] ), .B0(n2904), .Y(n2909)
         );
  OAI21X1 U2984 ( .A0(\decoder/w_PM_4[6] ), .A1(n2895), .B0(n2894), .Y(n2896)
         );
  AND2X2 U2986 ( .A(n669), .B(n2869), .Y(n1558) );
  AOI31X1 U2987 ( .A0(n2851), .A1(n695), .A2(n2850), .B0(n2849), .Y(n2854) );
  NAND3XL U2988 ( .A(n2846), .B(n709), .C(n2845), .Y(n2847) );
  OA22X2 U2989 ( .A0(\decoder/w_PM_1[5] ), .A1(n2835), .B0(n2872), .B1(
        \decoder/w_PM_1[6] ), .Y(n2846) );
  OAI22X1 U2990 ( .A0(\decoder/w_PM_1[3] ), .A1(n2869), .B0(n2834), .B1(n711), 
        .Y(n2839) );
  AOI21X1 U2991 ( .A0(n2869), .A1(\decoder/w_PM_1[3] ), .B0(n2833), .Y(n2840)
         );
  OAI21X1 U2992 ( .A0(\decoder/w_PM_2[6] ), .A1(n2904), .B0(n2866), .Y(n2860)
         );
  AOI21X1 U2993 ( .A0(n695), .A1(n2851), .B0(n2849), .Y(n2829) );
  MXI2X1 U2995 ( .A(n1084), .B(n1086), .S0(n1102), .Y(n699) );
  OAI21X1 U2996 ( .A0(n696), .A1(n2823), .B0(n2850), .Y(n2826) );
  OAI211XL U2997 ( .A0(n2824), .A1(n711), .B0(n2809), .C0(n2808), .Y(n2810) );
  MXI2X1 U2998 ( .A(n1416), .B(n1414), .S0(n1100), .Y(n686) );
  AND3X2 U2999 ( .A(n2805), .B(n682), .C(n2804), .Y(n2815) );
  OAI21X1 U3008 ( .A0(n3067), .A1(\decoder/u_ACS_matrix/w_PM_7_to_8_1[0] ), 
        .B0(n2486), .Y(n2524) );
  AOI21X1 U3009 ( .A0(n2482), .A1(n2485), .B0(n2496), .Y(n2497) );
  BUFX2 U3010 ( .A(n2432), .Y(n1204) );
  OAI21X1 U3013 ( .A0(n1937), .A1(\decoder/u_ACS_matrix/w_PM_4_to_5_4[2] ), 
        .B0(n1936), .Y(n1982) );
  OAI21X1 U3017 ( .A0(n2272), .A1(\decoder/u_ACS_matrix/w_PM_5_to_6_1[3] ), 
        .B0(n2284), .Y(n2317) );
  AOI21X1 U3018 ( .A0(n2269), .A1(n2276), .B0(n2315), .Y(n2282) );
  AOI21X1 U3023 ( .A0(n2648), .A1(n2647), .B0(n2615), .Y(n2616) );
  BUFX2 U3024 ( .A(n2599), .Y(n1228) );
  MX2X1 U3025 ( .A(n1534), .B(n1532), .S0(n1530), .Y(n1162) );
  MX2X1 U3026 ( .A(n1448), .B(n1450), .S0(n1460), .Y(n1166) );
  MX2X1 U3027 ( .A(n1456), .B(n1458), .S0(n1460), .Y(n1167) );
  MX2X1 U3028 ( .A(n1442), .B(n1444), .S0(n1460), .Y(n1168) );
  MX2X1 U3029 ( .A(n1452), .B(n1454), .S0(n1460), .Y(n1169) );
  MX2X1 U3030 ( .A(n1387), .B(n1385), .S0(n1327), .Y(n1170) );
  MX2X1 U3031 ( .A(n1408), .B(n1406), .S0(n1327), .Y(n1171) );
  MX2X1 U3032 ( .A(n1420), .B(n1418), .S0(n1327), .Y(n1172) );
  MX2X1 U3033 ( .A(n1094), .B(n1097), .S0(n978), .Y(n1173) );
  MX2X1 U3034 ( .A(n1432), .B(n1430), .S0(n978), .Y(n1175) );
  MX2X1 U3035 ( .A(n1456), .B(n1458), .S0(n2974), .Y(n1176) );
  MX2X1 U3036 ( .A(n1442), .B(n1444), .S0(n2974), .Y(n1178) );
  MX2X1 U3037 ( .A(n1448), .B(n1450), .S0(n2974), .Y(n1179) );
  MX2X1 U3038 ( .A(n1452), .B(n1454), .S0(n2974), .Y(n1180) );
  AND2X2 U3039 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_3[3] ), .B(
        \decoder/u_ACS_matrix/w_PM_5_to_6_3[4] ), .Y(n1184) );
  BUFX2 U3040 ( .A(n2595), .Y(n1229) );
  MXI2X1 U3044 ( .A(n1323), .B(n1325), .S0(n3007), .Y(n704) );
  AND3X2 U3062 ( .A(n2882), .B(n682), .C(n2881), .Y(n2822) );
  MXI2X1 U3089 ( .A(n1412), .B(n1410), .S0(n3007), .Y(n701) );
  OAI21X1 U3102 ( .A0(n682), .A1(n2863), .B0(n2884), .Y(n2876) );
  MXI2X1 U3106 ( .A(n1515), .B(n1513), .S0(n3007), .Y(n702) );
  MXI2X1 U3116 ( .A(n1466), .B(n1464), .S0(n3007), .Y(n703) );
  MXI2X1 U3132 ( .A(n1488), .B(n1486), .S0(n3007), .Y(n700) );
  AOI21X1 U3177 ( .A0(n2870), .A1(n669), .B0(n2869), .Y(n2873) );
  OAI2B1X1 U3198 ( .A1N(n1612), .A0(n975), .B0(n1810), .Y(n1600) );
  MXI2X1 U3200 ( .A(n2412), .B(n1147), .S0(n1120), .Y(n763) );
  AND2X2 U3204 ( .A(n2101), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[1] ), .Y(
        n1604) );
  OAI22X1 U3205 ( .A0(n1783), .A1(n1763), .B0(n1786), .B1(n1754), .Y(n926) );
  MXI2X1 U3206 ( .A(n1788), .B(n1787), .S0(n1786), .Y(n928) );
  MXI2X1 U3209 ( .A(n1787), .B(n1788), .S0(n1730), .Y(n911) );
  MXI2X1 U3210 ( .A(n1719), .B(n1726), .S0(n1730), .Y(n909) );
  MXI2X1 U3213 ( .A(n1798), .B(n971), .S0(n1793), .Y(n919) );
  MXI2X1 U3214 ( .A(n1796), .B(n1795), .S0(n1793), .Y(n918) );
  MXI2X1 U3216 ( .A(n1725), .B(n1724), .S0(n2919), .Y(n901) );
  NOR2BX1 U3217 ( .AN(\decoder/u_ACS_matrix/w_data_3_to_4_4[1] ), .B(n2936), 
        .Y(n885) );
  NOR2BX1 U3221 ( .AN(n2521), .B(n2520), .Y(n680) );
  MXI2X1 U3228 ( .A(n1728), .B(n1727), .S0(n1730), .Y(n910) );
  ACHCINX2 U3229 ( .CIN(n1814), .A(n1819), .B(n1822), .CO(n1815) );
  DFFSQXL R_251 ( .D(n2970), .CK(io_clk), .SN(n1634), .Q(n1323) );
  DFFSQXL R_170 ( .D(n2942), .CK(io_clk), .SN(n1634), .Q(n1420) );
  DFFSQXL R_69 ( .D(n1913), .CK(io_clk), .SN(n1634), .Q(n1534) );
  DFFSQXL R_70 ( .D(n1912), .CK(io_clk), .SN(n1634), .Q(n1532) );
  DFFSQXL R_250 ( .D(n2971), .CK(io_clk), .SN(n1631), .Q(n1325) );
  DFFSQXL R_171 ( .D(n2941), .CK(io_clk), .SN(n1635), .Q(n1418) );
  DFFSQXL R_183 ( .D(n2925), .CK(io_clk), .SN(n1635), .Q(n1406) );
  DFFSQXL R_200 ( .D(n2248), .CK(io_clk), .SN(n1634), .Q(n1385) );
  DFFSQXL R_182 ( .D(n2926), .CK(io_clk), .SN(n1635), .Q(n1408) );
  DFFSQXL R_168 ( .D(n2966), .CK(io_clk), .SN(n1632), .Q(n1422) );
  DFFSQXL R_207 ( .D(n2929), .CK(io_clk), .SN(n1635), .Q(n1373) );
  DFFSQXL R_205 ( .D(n2792), .CK(io_clk), .SN(n1634), .Q(n1377) );
  DFFSQXL R_149 ( .D(n2958), .CK(io_clk), .SN(n1635), .Q(n1456) );
  DFFSQXL R_151 ( .D(n2947), .CK(io_clk), .SN(n1635), .Q(n1452) );
  DFFSQXL R_153 ( .D(n2931), .CK(io_clk), .SN(n1634), .Q(n1448) );
  DFFSQXL R_156 ( .D(n2794), .CK(io_clk), .SN(n1635), .Q(n1442) );
  DFFSQXL R_199 ( .D(n2249), .CK(io_clk), .SN(n1634), .Q(n1387) );
  DFFSQXL R_148 ( .D(n2957), .CK(io_clk), .SN(n1635), .Q(n1458) );
  DFFSQXL R_155 ( .D(n2793), .CK(io_clk), .SN(n1634), .Q(n1444) );
  DFFSQXL R_53 ( .D(n2967), .CK(io_clk), .SN(n1635), .Q(n1546) );
  DFFSQXL R_152 ( .D(n2930), .CK(io_clk), .SN(n1635), .Q(n1450) );
  DFFSQXL R_150 ( .D(n2946), .CK(io_clk), .SN(n1634), .Q(n1454) );
  DFFSQXL R_90 ( .D(n2949), .CK(io_clk), .SN(n1634), .Q(n1513) );
  DFFSQXL R_118 ( .D(n2798), .CK(io_clk), .SN(n1634), .Q(n1486) );
  DFFSQXL R_139 ( .D(n2961), .CK(io_clk), .SN(n1634), .Q(n1464) );
  DFFSQXL R_180 ( .D(n2933), .CK(io_clk), .SN(n1635), .Q(n1410) );
  DFFSQXL R_209 ( .D(n2945), .CK(io_clk), .SN(n1635), .Q(n1369) );
  DFFSQXL R_211 ( .D(n2956), .CK(io_clk), .SN(n1634), .Q(n1365) );
  DFFSQXL R_162 ( .D(n1889), .CK(io_clk), .SN(n1635), .Q(n1430) );
  DFFSQXL R_161 ( .D(n1890), .CK(io_clk), .SN(n1635), .Q(n1432) );
  OAI2B1X2 U1602 ( .A1N(n2722), .A0(\decoder/u_ACS_matrix/w_PM_7_to_8_3[0] ), 
        .B0(n2713), .Y(n2787) );
  NAND3X4 U2324 ( .A(n1254), .B(n1253), .C(n2755), .Y(n1252) );
  INVX4 U1350 ( .A(n1252), .Y(n2771) );
  SDFFRHQX8 R_255 ( .D(\decoder/u_input_shifter/U_input_split/N51 ), .SI(1'b0), 
        .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(\decoder/w_enc_bit_8[0] ) );
  NAND3X2 U1685 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_3[0] ), .B(n2720), .C(
        n2723), .Y(n2726) );
  MXI2XL U2861 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_3[3] ), .B(n1213), 
        .S0(n2981), .Y(n1222) );
  MXI2XL U2862 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_3[4] ), .B(n1214), 
        .S0(n2981), .Y(n1223) );
  MXI2XL U2863 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_3[5] ), .B(n1212), 
        .S0(n2981), .Y(n1221) );
  MXI2XL U2874 ( .A(\decoder/u_ACS_matrix/w_data_7_to_8_3[6] ), .B(n1215), 
        .S0(n2981), .Y(n1224) );
  INVX3 U2092 ( .A(n1298), .Y(n1217) );
  SDFFSHQX4 R_30 ( .D(n3030), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1626), 
        .Q(n1561) );
  SDFFSHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_4/u_MEM/data_out_reg[7]  ( 
        .D(n1224), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1625), .Q(n993) );
  SDFFSHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_4/u_MEM/data_out_reg[6]  ( 
        .D(n1221), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1633), .Q(n3078) );
  SDFFSHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_4/u_MEM/data_out_reg[5]  ( 
        .D(n1223), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), .Q(n3076) );
  SDFFSHQX2 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_4/u_MEM/data_out_reg[4]  ( 
        .D(n1222), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), .Q(n3074) );
  SDFFRHQX2 \decoder/u_cmp_sel/data_out_reg[1]  ( .D(\decoder/u_cmp_sel/N43 ), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .Q(io_data_dec[1]) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/PM_out_reg[0]  ( 
        .D(n788), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_3[0] ) );
  OAI21X4 U2100 ( .A0(n2727), .A1(\decoder/u_ACS_matrix/w_PM_7_to_8_4[3] ), 
        .B0(n2731), .Y(n2779) );
  NAND3X4 U2422 ( .A(n2729), .B(n2730), .C(n2728), .Y(n2781) );
  NAND2BX4 U2452 ( .AN(n2662), .B(n2665), .Y(n2707) );
  INVX2 U1777 ( .A(n2727), .Y(n2729) );
  NAND2X2 U2412 ( .A(n2750), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_4[5] ), .Y(
        n2751) );
  OAI21X6 U1592 ( .A0(n2679), .A1(n1055), .B0(
        \decoder/u_ACS_matrix/w_PM_7_to_8_4[6] ), .Y(n1056) );
  CLKNAND2X2 U2413 ( .A(n2759), .B(n2758), .Y(n1253) );
  NOR2X8 U2148 ( .A(n994), .B(n2549), .Y(n2188) );
  CLKINVX2 U2101 ( .A(n1300), .Y(n1218) );
  OAI31X4 U1593 ( .A0(n2679), .A1(\decoder/u_ACS_matrix/w_PM_7_to_8_4[6] ), 
        .A2(n1055), .B0(n1056), .Y(n2688) );
  SDFFRQX4 \decoder/u_ACS_matrix/u_ACS_col_8/u_ACS_mem_1/u_MEM/data_out_reg[2]  ( 
        .D(n719), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/w_data_1[2] ) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_4/u_MEM/PM_out_reg[3]  ( 
        .D(n723), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_4[3] ) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/PM_out_reg[2]  ( 
        .D(n774), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_4[2] ) );
  SDFFSX1 R_179 ( .D(n1166), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1627), 
        .Q(n1412) );
  SDFFSX1 R_138 ( .D(n1167), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1629), 
        .Q(n1466) );
  SDFFSX1 R_117 ( .D(n1168), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1628), 
        .Q(n1488) );
  SDFFSX1 R_89 ( .D(n1169), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1626), .Q(
        n1515) );
  SDFFSX1 R_167 ( .D(n1182), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1630), 
        .Q(n1424) );
  SDFFSX1 R_210 ( .D(n1176), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1626), 
        .Q(n1367) );
  SDFFSX1 R_208 ( .D(n1180), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1371) );
  SDFFSX1 R_206 ( .D(n1179), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1629), 
        .Q(n1375) );
  SDFFSX1 R_204 ( .D(n1178), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1379) );
  SDFFSX1 R_288 ( .D(n2938), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1625), 
        .Q(n1094) );
  SDFFRX1 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_4/u_MEM/data_out_reg[1]  ( 
        .D(n1462), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1625), .QN(n2967)
         );
  SDFFRX1 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_4/u_MEM/data_out_reg[1]  ( 
        .D(n1462), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_4[1] ) );
  SDFFRX1 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_2/u_MEM/data_out_reg[1]  ( 
        .D(n1462), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_2[1] ) );
  SDFFRX1 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_2/u_MEM/data_out_reg[1]  ( 
        .D(n1462), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .QN(n2939)
         );
  SDFFRX1 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_2/u_MEM/data_out_reg[1]  ( 
        .D(n1462), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_data_3_to_4_2[1] ) );
  SDFFRX1 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_4/u_MEM/data_out_reg[1]  ( 
        .D(n1462), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_data_3_to_4_4[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/PM_out_reg[6]  ( 
        .D(n733), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n3039), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[6] ) );
  SDFFSX4 R_296 ( .D(
        \decoder/u_ACS_matrix/u_ACS_col_1/u_ACS_mem_3/u_ACS/ham_dist_2[0] ), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n3039), .QN(
        \decoder/u_ACS_matrix/w_PM_1_to_2_4[0] ) );
  SDFFSX1 R_154 ( .D(n2981), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1631), 
        .Q(n3032) );
  SDFFSHQX8 R_28 ( .D(n1127), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1631), 
        .Q(n1565) );
  SDFFSQX1 R_43 ( .D(n2378), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1550) );
  SDFFSHQX8 R_235 ( .D(n2964), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1338) );
  SDFFSHQX1 R_239 ( .D(n2384), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1629), 
        .Q(n1332) );
  SDFFSHQX8 R_92 ( .D(n1005), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1511) );
  NAND2BX8 U1877 ( .AN(n2546), .B(n1129), .Y(n2174) );
  MXI2X6 U1672 ( .A(n1525), .B(n1523), .S0(n1521), .Y(n796) );
  NAND2X4 U2605 ( .A(n1024), .B(n2342), .Y(n2339) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_2/u_MEM/PM_out_reg[0]  ( 
        .D(n843), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_2[0] ) );
  NAND2X6 U1865 ( .A(n2188), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[3] ), .Y(
        n2190) );
  INVX2 U2062 ( .A(n669), .Y(n2891) );
  NAND2X2 U2186 ( .A(n2724), .B(n2723), .Y(n2725) );
  INVX4 U2456 ( .A(n3067), .Y(n2720) );
  AOI2BB2X4 U1849 ( .B0(n1121), .B1(n671), .A0N(n2890), .A1N(n697), .Y(n1125)
         );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_3/u_MEM/PM_out_reg[1]  ( 
        .D(n787), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_3[1] ) );
  SDFFSHQX4 R_213 ( .D(n2516), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1361) );
  SDFFSHQX4 R_136 ( .D(n2535), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1468) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/PM_out_reg[2]  ( 
        .D(n809), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_1[2] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/data_out_reg[2]  ( 
        .D(n769), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1635), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_1[2] ) );
  SDFFSHQX2 R_142 ( .D(n1127), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1460) );
  SDFFSHQX4 R_128 ( .D(n1127), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1632), 
        .Q(n1476) );
  SDFFSQX2 R_297 ( .D(n2920), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1634), 
        .Q(n1076) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_4/u_MEM/PM_out_reg[0]  ( 
        .D(n822), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_1/u_MEM/PM_out_reg[2]  ( 
        .D(n926), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_1[2] ) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_4/u_MEM/PM_out_reg[2]  ( 
        .D(n862), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_4_to_5_4[2] ) );
  SDFFRQX4 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_3/u_MEM/data_out_reg[2]  ( 
        .D(n836), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_data_5_to_6_3[2] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_4/u_ACS_mem_4/u_MEM/data_out_reg[2]  ( 
        .D(n1191), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_data_4_to_5_4[2] ) );
  SDFFRHQX2 \decoder/u_cmp_sel/data_out_reg[3]  ( .D(\decoder/u_cmp_sel/N45 ), 
        .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(io_data_dec[3]) );
  SDFFSHQX8 R_289 ( .D(n2999), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1625), 
        .Q(n1092) );
  NOR2X2 U2877 ( .A(n1148), .B(n1174), .Y(n2770) );
  MXI2X8 U1670 ( .A(n1502), .B(n1500), .S0(n1498), .Y(n797) );
  XNOR2X4 U2098 ( .A(n2751), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_4[6] ), .Y(
        n2765) );
  INVX3 U2424 ( .A(n2737), .Y(n1299) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/PM_out_reg[0]  ( 
        .D(n764), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[0] ) );
  NAND3X2 U1098 ( .A(n1027), .B(n2747), .C(n2746), .Y(n2758) );
  INVX4 U1099 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_1[0] ), .Y(n2988) );
  AOI2B1X2 U1100 ( .A1N(n2988), .A0(n2473), .B0(n2488), .Y(n2428) );
  INVX2 U1105 ( .A(n1174), .Y(n2990) );
  AND2X6 U1108 ( .A(n2763), .B(n2990), .Y(n2767) );
  AO21X4 U1109 ( .A0(n1803), .A1(n1804), .B0(n1891), .Y(n2991) );
  OAI21X4 U1114 ( .A0(n1892), .A1(\decoder/u_ACS_matrix/w_PM_3_to_4_2[1] ), 
        .B0(n1909), .Y(n1919) );
  MXI2X2 U1117 ( .A(n2089), .B(n2088), .S0(n2952), .Y(n822) );
  CLKNAND2X4 U1118 ( .A(n1964), .B(n1966), .Y(n1846) );
  OAI21XL U1121 ( .A0(n1802), .A1(\decoder/u_ACS_matrix/w_PM_3_to_4_2[1] ), 
        .B0(n1813), .Y(n2992) );
  OAI21X1 U1122 ( .A0(n1802), .A1(\decoder/u_ACS_matrix/w_PM_3_to_4_2[1] ), 
        .B0(n1813), .Y(n1823) );
  INVX2 U1126 ( .A(n1823), .Y(n1807) );
  OAI21X3 U1132 ( .A0(n1910), .A1(n1914), .B0(n1917), .Y(n1916) );
  AOI21X4 U1135 ( .A0(n1905), .A1(n1904), .B0(n1907), .Y(n1914) );
  CLKAND2X4 U1137 ( .A(n1801), .B(n1185), .Y(n1818) );
  MXI2X8 U1139 ( .A(n1404), .B(n1402), .S0(n1092), .Y(n863) );
  OAI21X2 U1143 ( .A0(n1899), .A1(\decoder/u_ACS_matrix/w_PM_3_to_4_1[1] ), 
        .B0(n1904), .Y(n1918) );
  NAND2X4 U1152 ( .A(n1899), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_1[1] ), .Y(
        n1904) );
  CLKAND2X2 U1153 ( .A(n2920), .B(\decoder/u_ACS_matrix/w_data_3_to_4_2[1] ), 
        .Y(n895) );
  INVXL U1154 ( .A(n1807), .Y(n1134) );
  NAND2X6 U1162 ( .A(n2012), .B(n2011), .Y(n2993) );
  MXI2XL U1163 ( .A(n2099), .B(n2063), .S0(n2098), .Y(n839) );
  OAI2B1X4 U1164 ( .A1N(n1612), .A0(n975), .B0(n1810), .Y(n1824) );
  BUFX3 U1166 ( .A(n1801), .Y(n975) );
  NAND2X2 U1168 ( .A(n1801), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_1[1] ), .Y(
        n1810) );
  NOR2X6 U1170 ( .A(n1813), .B(n1908), .Y(n1812) );
  NAND2X8 U1174 ( .A(n2102), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[3] ), .Y(
        n2127) );
  NAND2BX8 U1175 ( .AN(n1818), .B(n1811), .Y(n1819) );
  NOR2X4 U1182 ( .A(n2127), .B(n2285), .Y(n2166) );
  NOR2X2 U1196 ( .A(n2157), .B(n2159), .Y(n2113) );
  NOR2BX2 U1201 ( .AN(n1824), .B(n2992), .Y(n1809) );
  AOI21X3 U1203 ( .A0(n2994), .A1(n1813), .B0(n1812), .Y(n1822) );
  CLKINVX40 U1204 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_2[2] ), .Y(n2994) );
  CLKNAND2X4 U1205 ( .A(n2156), .B(n2123), .Y(n2124) );
  OAI21X4 U1206 ( .A0(n2164), .A1(n2165), .B0(n2163), .Y(n2008) );
  OAI21X4 U1210 ( .A0(n1991), .A1(\decoder/u_ACS_matrix/w_PM_5_to_6_3[3] ), 
        .B0(n2007), .Y(n2146) );
  NAND2BX8 U1211 ( .AN(n2166), .B(n2118), .Y(n2150) );
  INVX1 U1216 ( .A(n2150), .Y(n2154) );
  OR2X4 U1224 ( .A(n1992), .B(n1274), .Y(n2995) );
  NAND2X3 U1234 ( .A(n1997), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_4[1] ), .Y(
        n1992) );
  INVXL U1235 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_4[2] ), .Y(n1274) );
  OAI2BB1X2 U1248 ( .A0N(n2156), .A1N(n3089), .B0(n2155), .Y(n784) );
  OAI21X4 U1251 ( .A0(n2162), .A1(n2160), .B0(n2161), .Y(n2009) );
  OAI21X2 U1253 ( .A0(n2102), .A1(\decoder/u_ACS_matrix/w_PM_5_to_6_1[3] ), 
        .B0(n2127), .Y(n2159) );
  NOR2X8 U1255 ( .A(n2105), .B(n2270), .Y(n2102) );
  OAI21X1 U1263 ( .A0(n2226), .A1(n3001), .B0(n2311), .Y(n2227) );
  CLKINVX4 U1265 ( .A(n2215), .Y(n2327) );
  INVX3 U1267 ( .A(n2550), .Y(n2564) );
  AND2X1 U1268 ( .A(n2571), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_4[5] ), .Y(
        n1072) );
  INVX8 U1270 ( .A(n2385), .Y(n2176) );
  NAND2BX1 U1275 ( .AN(n695), .B(n668), .Y(n2879) );
  INVX4 U1283 ( .A(n1118), .Y(n991) );
  INVX4 U1284 ( .A(n991), .Y(n992) );
  NAND2X1 U1286 ( .A(n2653), .B(n2573), .Y(n2572) );
  MXI2XL U1287 ( .A(n2319), .B(n2318), .S0(n2955), .Y(n809) );
  NAND3X4 U1296 ( .A(n1199), .B(n2560), .C(n2559), .Y(n2562) );
  NAND2BX4 U1297 ( .AN(n2578), .B(n2577), .Y(n1199) );
  MXI2X1 U1306 ( .A(n2580), .B(n3098), .S0(n2400), .Y(n751) );
  AOI21XL U1307 ( .A0(n1713), .A1(n1712), .B0(n1711), .Y(n1729) );
  OAI21X1 U1312 ( .A0(n2076), .A1(n2016), .B0(n2015), .Y(n2038) );
  OAI21X2 U1314 ( .A0(n1610), .A1(\decoder/u_ACS_matrix/w_PM_4_to_5_2[3] ), 
        .B0(n2077), .Y(n2081) );
  MXI2XL U1315 ( .A(n2991), .B(n1920), .S0(n1132), .Y(n874) );
  NOR2BX4 U1318 ( .AN(n1782), .B(n1781), .Y(n1783) );
  BUFX2 U1319 ( .A(n2067), .Y(n2996) );
  AOI21XL U1320 ( .A0(n1933), .A1(n1976), .B0(n1952), .Y(n818) );
  CLKINVX2 U1321 ( .A(n1861), .Y(n1957) );
  OAI211X4 U1324 ( .A0(n1761), .A1(n1751), .B0(n1714), .C0(n1758), .Y(n1718)
         );
  NAND2BX4 U1327 ( .AN(n1727), .B(n1728), .Y(n1714) );
  MXI2XL U1328 ( .A(n1163), .B(n1906), .S0(n1132), .Y(n871) );
  NOR2X3 U1329 ( .A(n1938), .B(n1133), .Y(n1935) );
  CLKAND2X4 U1331 ( .A(n2937), .B(\decoder/u_ACS_matrix/w_data_3_to_4_4[1] ), 
        .Y(n1191) );
  CLKINVX4 U1335 ( .A(n890), .Y(n2014) );
  AOI21XL U1348 ( .A0(n1620), .A1(n1988), .B0(n2165), .Y(n771) );
  INVXL U1349 ( .A(n2061), .Y(n2997) );
  INVX2 U1355 ( .A(n2096), .Y(n2061) );
  OAI21X4 U1357 ( .A0(n2058), .A1(n861), .B0(n2063), .Y(n2096) );
  NOR2X1 U1363 ( .A(n1983), .B(n1984), .Y(n1940) );
  MXI2XL U1367 ( .A(n1785), .B(n1784), .S0(n1786), .Y(n927) );
  AOI2B1X4 U1369 ( .A1N(n2048), .A0(n1133), .B0(n2056), .Y(n2090) );
  INVXL U1370 ( .A(n1903), .Y(n2998) );
  NAND2X4 U1371 ( .A(n2061), .B(n1154), .Y(n2072) );
  OAI21XL U1375 ( .A0(n1910), .A1(n1914), .B0(n1917), .Y(n982) );
  INVX3 U1377 ( .A(n1876), .Y(n1925) );
  OAI21X3 U1385 ( .A0(n2045), .A1(\decoder/u_ACS_matrix/w_PM_4_to_5_4[2] ), 
        .B0(n2057), .Y(n2092) );
  NAND2X4 U1386 ( .A(n2045), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_4[2] ), .Y(
        n2057) );
  INVX3 U1393 ( .A(n2049), .Y(n2045) );
  AOI2BB1X2 U1404 ( .A0N(n2993), .A1N(\decoder/u_ACS_matrix/w_PM_4_to_5_4[0] ), 
        .B0(n2044), .Y(n1946) );
  NOR2X1 U1410 ( .A(n1133), .B(n1938), .Y(n966) );
  OAI211X1 U1412 ( .A0(n1952), .A1(n1949), .B0(n1948), .C0(n1947), .Y(n1950)
         );
  NAND2X4 U1414 ( .A(n891), .B(n2024), .Y(n2019) );
  CLKINVX3 U1423 ( .A(n1924), .Y(n2999) );
  INVX3 U1440 ( .A(n1924), .Y(n2937) );
  MXI2XL U1444 ( .A(n1930), .B(n1929), .S0(n2999), .Y(n864) );
  CLKNAND2X2 U1451 ( .A(\decoder/w_enc_bit_4[0] ), .B(n1240), .Y(n1882) );
  NAND2BXL U1458 ( .AN(n1859), .B(n1975), .Y(n1321) );
  NAND2X4 U1461 ( .A(n1595), .B(n1596), .Y(n1859) );
  OAI21X8 U1462 ( .A0(n1903), .A1(n970), .B0(n1901), .Y(n1910) );
  INVX2 U1467 ( .A(n1919), .Y(n1903) );
  NAND2BX8 U1468 ( .AN(n1918), .B(n1900), .Y(n1901) );
  NAND3X3 U1469 ( .A(n1846), .B(n2023), .C(n2030), .Y(n1848) );
  NAND2X4 U1470 ( .A(n2022), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_2[1] ), .Y(
        n2021) );
  CLKINVX1 U1471 ( .A(n1137), .Y(n2029) );
  MXI2X1 U1474 ( .A(n2089), .B(n2088), .S0(n2953), .Y(n843) );
  MXI2XL U1476 ( .A(n1153), .B(n2091), .S0(n2953), .Y(n841) );
  MXI2XL U1479 ( .A(n2997), .B(n969), .S0(n2953), .Y(n840) );
  MXI2XL U1481 ( .A(n3000), .B(n2093), .S0(n2953), .Y(n842) );
  MXI2XL U1485 ( .A(n1175), .B(n1162), .S0(n2953), .Y(n844) );
  MXI2XL U1487 ( .A(n2924), .B(n2923), .S0(n2953), .Y(n845) );
  NAND3X3 U1493 ( .A(n2073), .B(n2062), .C(n2072), .Y(n2074) );
  BUFX2 U1498 ( .A(n2012), .Y(n1137) );
  AOI21X6 U1504 ( .A0(n2025), .A1(n1135), .B0(n2010), .Y(n2024) );
  AOI21X2 U1510 ( .A0(n2026), .A1(n2025), .B0(n986), .Y(n2033) );
  OAI21X2 U1512 ( .A0(n891), .A1(n1850), .B0(n1849), .Y(n1962) );
  NAND3X2 U1519 ( .A(n1852), .B(n1853), .C(n1855), .Y(n1857) );
  NAND2X8 U1522 ( .A(n1845), .B(\decoder/u_ACS_matrix/w_PM_4_to_5_1[0] ), .Y(
        n2025) );
  MXI2XL U1524 ( .A(n1961), .B(n1960), .S0(n1958), .Y(n830) );
  NAND2X3 U1525 ( .A(n1959), .B(n1961), .Y(n1855) );
  MXI2XL U1532 ( .A(n2998), .B(n1918), .S0(n1132), .Y(n873) );
  NAND2BX8 U1534 ( .AN(n1919), .B(n1902), .Y(n1900) );
  MXI2XL U1535 ( .A(n1966), .B(n1965), .S0(n1958), .Y(n832) );
  INVXL U1550 ( .A(n1133), .Y(n968) );
  MXI2XL U1551 ( .A(n1979), .B(n1978), .S0(n2952), .Y(n819) );
  MXI2XL U1559 ( .A(n2924), .B(n2923), .S0(n2952), .Y(n824) );
  MXI2XL U1565 ( .A(n1175), .B(n1162), .S0(n2952), .Y(n823) );
  MXI2XL U1574 ( .A(n1985), .B(n1984), .S0(n2952), .Y(n821) );
  MXI2XL U1577 ( .A(n1141), .B(n1981), .S0(n2952), .Y(n820) );
  MXI2XL U1580 ( .A(n2041), .B(n2040), .S0(n1958), .Y(n834) );
  XNOR2X4 U1585 ( .A(n1849), .B(n890), .Y(n1959) );
  INVXL U1587 ( .A(n2053), .Y(n3000) );
  OAI31X1 U1589 ( .A0(n2066), .A1(n2044), .A2(n863), .B0(n1054), .Y(n2094) );
  NAND2X3 U1590 ( .A(n891), .B(n1850), .Y(n1849) );
  MXI2XL U1611 ( .A(n2922), .B(n2921), .S0(n1958), .Y(n835) );
  AOI2BB2X4 U1614 ( .B0(n2146), .B1(n1042), .A0N(n1028), .A1N(n2145), .Y(n773)
         );
  NOR2XL U1626 ( .A(n2940), .B(n2939), .Y(n857) );
  MXI2X1 U1627 ( .A(n2087), .B(n2086), .S0(n2940), .Y(n854) );
  NAND3BX4 U1638 ( .AN(n2035), .B(n2034), .C(n2037), .Y(n2036) );
  AOI21X2 U1641 ( .A0(n1844), .A1(n2025), .B0(n1850), .Y(n1964) );
  AOI21X3 U1643 ( .A0(n2025), .A1(n1137), .B0(n2010), .Y(n1850) );
  OAI21XL U1649 ( .A0(\decoder/u_ACS_matrix/w_PM_3_to_4_3[0] ), .A1(n1804), 
        .B0(n1863), .Y(n1930) );
  CLKNAND2X2 U1652 ( .A(n1863), .B(n1882), .Y(n1739) );
  INVX6 U1653 ( .A(n2050), .Y(n2044) );
  OAI21XL U1665 ( .A0(n2066), .A1(n2044), .B0(n981), .Y(n1054) );
  XNOR2XL U1667 ( .A(n1997), .B(n2220), .Y(n2141) );
  INVXL U1668 ( .A(n2157), .Y(n2158) );
  XNOR2X4 U1673 ( .A(n1604), .B(n2270), .Y(n2147) );
  CLKNAND2X2 U1683 ( .A(n2090), .B(n2092), .Y(n2068) );
  AOI2B1XL U1693 ( .A1N(\decoder/u_ACS_matrix/w_PM_3_to_4_1[0] ), .A0(n1804), 
        .B0(n3091), .Y(n1049) );
  MXI2XL U1694 ( .A(n1912), .B(n1913), .S0(n2920), .Y(n894) );
  MXI2XL U1697 ( .A(n1920), .B(n2991), .S0(n2920), .Y(n893) );
  MXI2XL U1711 ( .A(n1600), .B(n1134), .S0(n2920), .Y(n892) );
  NAND2BX1 U1725 ( .AN(n2079), .B(n2078), .Y(n2080) );
  NAND2X4 U1733 ( .A(n1184), .B(n2212), .Y(n2328) );
  CLKNAND2X2 U1734 ( .A(n2239), .B(n2216), .Y(n2247) );
  NAND2X4 U1737 ( .A(n1802), .B(\decoder/u_ACS_matrix/w_PM_3_to_4_2[1] ), .Y(
        n1813) );
  OAI22X2 U1738 ( .A0(n1809), .A1(n1808), .B0(n1807), .B1(n1600), .Y(n1814) );
  MXI2XL U1749 ( .A(n2922), .B(n2921), .S0(n2940), .Y(n856) );
  MXI2XL U1751 ( .A(n2041), .B(n2040), .S0(n2940), .Y(n855) );
  MXI2XL U1752 ( .A(n2077), .B(n2076), .S0(n2940), .Y(n850) );
  MXI2XL U1761 ( .A(n2083), .B(n2082), .S0(n2940), .Y(n852) );
  MXI2XL U1771 ( .A(n2085), .B(n2084), .S0(n2940), .Y(n853) );
  NOR2X1 U1807 ( .A(n2146), .B(n2145), .Y(n2004) );
  NAND2X3 U1825 ( .A(n2008), .B(n2161), .Y(n1308) );
  INVXL U1843 ( .A(n2228), .Y(n3001) );
  CLKNAND2X2 U1853 ( .A(n2120), .B(n2119), .Y(n2122) );
  NOR2X2 U1859 ( .A(n2148), .B(n2147), .Y(n2104) );
  BUFX2 U1866 ( .A(n2148), .Y(n1149) );
  CLKNAND2X2 U1867 ( .A(n2147), .B(n2148), .Y(n2112) );
  XNOR2X4 U1872 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_3[4] ), .B(n2237), .Y(
        n2300) );
  NAND2BX1 U1878 ( .AN(n2326), .B(n2240), .Y(n2243) );
  NAND2BX2 U1884 ( .AN(n2308), .B(n2230), .Y(n2229) );
  BUFX6 U1885 ( .A(n2024), .Y(n986) );
  AOI21X4 U1890 ( .A0(n2019), .A1(n2014), .B0(n2039), .Y(n2078) );
  INVX3 U1891 ( .A(n2039), .Y(n2076) );
  NOR2X4 U1892 ( .A(n2014), .B(n2019), .Y(n2039) );
  MXI2XL U1893 ( .A(n2576), .B(n2575), .S0(n1127), .Y(n722) );
  OAI211X1 U1896 ( .A0(n2085), .A1(n2033), .B0(n2032), .C0(n2031), .Y(n1053)
         );
  MXI2XL U1898 ( .A(n1179), .B(n2929), .S0(n3092), .Y(n688) );
  MXI2XL U1900 ( .A(n1178), .B(n2792), .S0(n3092), .Y(n687) );
  MXI2XL U1902 ( .A(n1182), .B(n2966), .S0(n2977), .Y(n691) );
  MXI2XL U1907 ( .A(n1176), .B(n2956), .S0(n2977), .Y(n690) );
  MXI2XL U1911 ( .A(n1180), .B(n2945), .S0(n2977), .Y(n689) );
  NAND3X4 U1915 ( .A(n2515), .B(n2513), .C(n2514), .Y(n1126) );
  NAND2X4 U1917 ( .A(n2101), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[1] ), .Y(
        n2105) );
  NAND2X2 U1924 ( .A(n2219), .B(n2225), .Y(n2222) );
  MXI2XL U1926 ( .A(n2149), .B(n1149), .S0(n2954), .Y(n786) );
  MXI2XL U1927 ( .A(n2299), .B(n2298), .S0(n3089), .Y(n789) );
  MXI2XL U1928 ( .A(n2928), .B(n2927), .S0(n3089), .Y(n790) );
  MXI2XL U1929 ( .A(n2944), .B(n2943), .S0(n3089), .Y(n791) );
  MXI2XL U1931 ( .A(n2159), .B(n2158), .S0(n2954), .Y(n785) );
  MXI2XL U1935 ( .A(n2323), .B(n2322), .S0(n2954), .Y(n788) );
  MXI2XL U1937 ( .A(n2132), .B(n2131), .S0(n2954), .Y(n787) );
  NAND2X3 U1942 ( .A(n2252), .B(n1314), .Y(n2101) );
  NOR3X2 U1945 ( .A(n2691), .B(n2692), .C(n2698), .Y(n2686) );
  BUFX6 U1946 ( .A(n2244), .Y(n1230) );
  AOI21XL U1948 ( .A0(n2226), .A1(n2209), .B0(n2311), .Y(n1996) );
  OAI21X2 U1949 ( .A0(n2310), .A1(n2228), .B0(n2227), .Y(n2230) );
  CLKNAND2X2 U1965 ( .A(n2225), .B(n2219), .Y(n1313) );
  CLKINVX2 U1967 ( .A(n776), .Y(n1557) );
  OAI21X4 U1968 ( .A0(n1124), .A1(n1144), .B0(n1307), .Y(n2536) );
  OAI21X2 U1978 ( .A0(n2496), .A1(\decoder/u_ACS_matrix/w_PM_7_to_8_1[3] ), 
        .B0(n1310), .Y(n2535) );
  INVX3 U1986 ( .A(n670), .Y(n2890) );
  NOR2X8 U1987 ( .A(n2916), .B(n1145), .Y(n2983) );
  NOR2X4 U2013 ( .A(n2563), .B(n2544), .Y(n2571) );
  MXI2XL U2016 ( .A(n2654), .B(n2653), .S0(n1127), .Y(n721) );
  BUFX3 U2019 ( .A(n2527), .Y(n1139) );
  MXI2XL U2022 ( .A(n2323), .B(n2322), .S0(n2955), .Y(n811) );
  AOI21X2 U2025 ( .A0(n2663), .A1(n3085), .B0(n988), .Y(n2662) );
  NAND2X3 U2028 ( .A(n2707), .B(n2706), .Y(n2681) );
  OAI21XL U2034 ( .A0(n2558), .A1(n2579), .B0(n2557), .Y(n2559) );
  INVXL U2036 ( .A(n2642), .Y(n3002) );
  INVX2 U2040 ( .A(n3002), .Y(n3003) );
  NOR2X4 U2046 ( .A(n2386), .B(n1251), .Y(n1302) );
  INVX2 U2050 ( .A(n2185), .Y(n2186) );
  CLKAND2X2 U2051 ( .A(n1620), .B(\decoder/u_ACS_matrix/w_data_5_to_6_4[1] ), 
        .Y(n780) );
  MXI2XL U2054 ( .A(n2248), .B(n2249), .S0(n1620), .Y(n777) );
  MXI2XL U2061 ( .A(n2925), .B(n2926), .S0(n1620), .Y(n778) );
  MXI2XL U2074 ( .A(n2941), .B(n2942), .S0(n1620), .Y(n779) );
  CLKINVX4 U2076 ( .A(n2480), .Y(n1124) );
  CLKINVX8 U2081 ( .A(n1303), .Y(n958) );
  AOI2B1X1 U2087 ( .A1N(\decoder/u_ACS_matrix/w_PM_6_to_7_4[4] ), .A0(n2563), 
        .B0(n2571), .Y(n2569) );
  NOR2X1 U2095 ( .A(n2518), .B(n2533), .Y(n2452) );
  NOR2BXL U2104 ( .AN(n2519), .B(n2518), .Y(n707) );
  NOR2X2 U2109 ( .A(n2518), .B(n2459), .Y(n2460) );
  NAND2X4 U2111 ( .A(n1295), .B(n1601), .Y(n1294) );
  INVX2 U2113 ( .A(n2384), .Y(n2189) );
  INVX10 U2131 ( .A(n2167), .Y(n2177) );
  MXI2XL U2132 ( .A(n2382), .B(n2381), .S0(n2400), .Y(n747) );
  MXI2XL U2140 ( .A(n2387), .B(n2386), .S0(n2400), .Y(n750) );
  MXI2XL U2143 ( .A(n2380), .B(n2379), .S0(n2400), .Y(n746) );
  NOR2X1 U2146 ( .A(n2643), .B(n2620), .Y(n2621) );
  NAND2BX4 U2149 ( .AN(n685), .B(n3020), .Y(n2817) );
  INVX4 U2152 ( .A(n1098), .Y(n685) );
  CLKNAND2X2 U2162 ( .A(n1145), .B(n3088), .Y(n3087) );
  OAI22X2 U2166 ( .A0(n667), .A1(n2799), .B0(\decoder/w_PM_4[6] ), .B1(n2906), 
        .Y(n2863) );
  INVX1 U2167 ( .A(n667), .Y(n1002) );
  NOR2X3 U2169 ( .A(n2203), .B(n2189), .Y(n1245) );
  INVX3 U2170 ( .A(n2617), .Y(n3014) );
  OAI21X4 U2178 ( .A0(n1072), .A1(n2652), .B0(n2574), .Y(n1275) );
  NOR3X2 U2190 ( .A(n2691), .B(n2690), .C(n2692), .Y(n2684) );
  MXI2XL U2203 ( .A(n2534), .B(n2533), .S0(n2710), .Y(n708) );
  MXI2XL U2215 ( .A(n2525), .B(n2524), .S0(n2710), .Y(n713) );
  MXI2XL U2217 ( .A(n3027), .B(n2538), .S0(n2710), .Y(n710) );
  MXI2XL U2221 ( .A(n997), .B(n2529), .S0(n2710), .Y(n712) );
  CLKNAND2X2 U2223 ( .A(n2446), .B(n2445), .Y(n2453) );
  INVXL U2227 ( .A(n3024), .Y(n3004) );
  INVX2 U2244 ( .A(n3004), .Y(n3005) );
  NAND3BX2 U2254 ( .AN(n1558), .B(n2865), .C(n1125), .Y(n2868) );
  INVX3 U2264 ( .A(n3024), .Y(n3006) );
  NAND2X3 U2265 ( .A(n2543), .B(n2435), .Y(n2443) );
  NAND2BX2 U2281 ( .AN(n2516), .B(n2517), .Y(n2503) );
  OAI21X3 U2288 ( .A0(n1597), .A1(\decoder/u_ACS_matrix/w_PM_7_to_8_1[4] ), 
        .B0(n2475), .Y(n2516) );
  BUFX4 U2313 ( .A(n2255), .Y(n1314) );
  NOR2X3 U2321 ( .A(n2362), .B(n1194), .Y(n960) );
  MXI2X1 U2331 ( .A(n2646), .B(n2645), .S0(n1623), .Y(n737) );
  NAND2BX1 U2386 ( .AN(n2646), .B(n2645), .Y(n2629) );
  OAI21X8 U2389 ( .A0(n1198), .A1(\decoder/u_ACS_matrix/w_PM_6_to_7_3[0] ), 
        .B0(n2545), .Y(n2579) );
  OAI22X2 U2394 ( .A0(n698), .A1(n2887), .B0(n2892), .B1(n697), .Y(n2842) );
  OAI21X1 U2410 ( .A0(n2690), .A1(n2698), .B0(n2689), .Y(n2695) );
  NAND2BXL U2417 ( .AN(n2488), .B(n2471), .Y(n1599) );
  NOR2X3 U2425 ( .A(n2185), .B(n1302), .Y(n2200) );
  AOI31X4 U2427 ( .A0(n2568), .A1(n2567), .A2(n1280), .B0(n1278), .Y(n1277) );
  NAND2BXL U2429 ( .AN(\decoder/w_PM_1[5] ), .B(n667), .Y(n2897) );
  NAND2BX2 U2431 ( .AN(n681), .B(n667), .Y(n2882) );
  NOR2BX4 U2432 ( .AN(n667), .B(\decoder/w_PM_2[5] ), .Y(n2903) );
  DLY1X1 U2434 ( .A(n724), .Y(n988) );
  NAND2X6 U2438 ( .A(n1249), .B(n1248), .Y(n3025) );
  NAND2X4 U2443 ( .A(n1249), .B(n1248), .Y(n2254) );
  INVX4 U2446 ( .A(n1205), .Y(n2734) );
  NAND2BX2 U2451 ( .AN(n2267), .B(n2258), .Y(n3024) );
  NAND2BX2 U2459 ( .AN(n670), .B(n697), .Y(n2870) );
  DLY1X1 U2474 ( .A(n1102), .Y(n3007) );
  OAI22X4 U2479 ( .A0(n672), .A1(n2886), .B0(n671), .B1(n2887), .Y(n2889) );
  AND2X8 U2481 ( .A(n749), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_2[1] ), .Y(
        n1257) );
  MXI2X6 U2484 ( .A(n1554), .B(n1552), .S0(n1082), .Y(n749) );
  INVXL U2488 ( .A(n2168), .Y(n3008) );
  NAND2XL U2501 ( .A(n3008), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_4[3] ), .Y(
        n2184) );
  NAND2X4 U2507 ( .A(n3009), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[0] ), .Y(
        n2713) );
  CLKINVX3 U2511 ( .A(n2722), .Y(n3009) );
  OAI21X4 U2517 ( .A0(n2365), .A1(\decoder/u_ACS_matrix/w_PM_6_to_7_1[3] ), 
        .B0(n2364), .Y(n2408) );
  BUFX2 U2529 ( .A(n2905), .Y(n3010) );
  CLKINVX2 U2550 ( .A(n2304), .Y(n3011) );
  OAI2B11X4 U2558 ( .A1N(n3011), .A0(n2244), .B0(n2303), .C0(n2245), .Y(n1227)
         );
  NAND2X2 U2560 ( .A(n3012), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_2[3] ), .Y(
        n2120) );
  XNOR2X4 U2561 ( .A(n3012), .B(n2286), .Y(n2157) );
  NAND3X4 U2562 ( .A(n3013), .B(n2426), .C(n2425), .Y(n2446) );
  NAND2X2 U2565 ( .A(n2537), .B(n2422), .Y(n3013) );
  NAND4X4 U2570 ( .A(n2612), .B(n3014), .C(n2610), .D(n2609), .Y(n2628) );
  CLKINVX1 U2571 ( .A(n3015), .Y(n3016) );
  NAND2BX2 U2576 ( .AN(n2525), .B(n2524), .Y(n3015) );
  OAI211X2 U2578 ( .A0(n2530), .A1(n2528), .B0(n3015), .C0(n2433), .Y(n2434)
         );
  NAND3BX4 U2587 ( .AN(n3016), .B(n2492), .C(n2490), .Y(n2494) );
  OR2X8 U2600 ( .A(n1241), .B(n3017), .Y(n2289) );
  NOR2X3 U2601 ( .A(n1241), .B(n2286), .Y(n3018) );
  NAND2BX8 U2606 ( .AN(n2286), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_2[4] ), 
        .Y(n3017) );
  INVX5 U2614 ( .A(n2313), .Y(n2291) );
  OAI21X8 U2615 ( .A0(\decoder/u_ACS_matrix/w_PM_5_to_6_2[4] ), .A1(n3018), 
        .B0(n2289), .Y(n2313) );
  NAND3X2 U2616 ( .A(n2454), .B(n2453), .C(n2711), .Y(n2464) );
  NOR2BX2 U2619 ( .AN(n2599), .B(n2332), .Y(n2333) );
  NAND2BX1 U2620 ( .AN(\decoder/u_ACS_matrix/w_PM_6_to_7_1[1] ), .B(n1155), 
        .Y(n2332) );
  NAND2X4 U2625 ( .A(n2713), .B(n2721), .Y(n2735) );
  OAI2BB1X4 U2628 ( .A0N(\decoder/u_ACS_matrix/w_PM_7_to_8_1[1] ), .A1N(n2488), 
        .B0(n2418), .Y(n2419) );
  NAND3X2 U2638 ( .A(n2473), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_1[1] ), .C(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[0] ), .Y(n2418) );
  CLKNAND2X2 U2641 ( .A(n2486), .B(n1019), .Y(n2474) );
  INVX4 U2671 ( .A(\decoder/w_enc_bit_8[0] ), .Y(n3065) );
  NAND2X3 U2672 ( .A(n2331), .B(n1239), .Y(n2362) );
  XNOR2X2 U2677 ( .A(n2340), .B(n2175), .Y(n2558) );
  NOR2BX2 U2693 ( .AN(n960), .B(n2593), .Y(n2353) );
  NOR2BXL U2718 ( .AN(n2688), .B(n2702), .Y(n693) );
  DLY1X1 U2739 ( .A(n2578), .Y(n3019) );
  NOR2X8 U2766 ( .A(n726), .B(n1299), .Y(n1298) );
  NAND2X3 U2772 ( .A(n1440), .B(n1438), .Y(n1434) );
  BUFX14 U2841 ( .A(n2604), .Y(n1155) );
  NAND2X3 U2845 ( .A(n2336), .B(n2362), .Y(n2410) );
  NAND2BX1 U2846 ( .AN(\decoder/u_ACS_matrix/w_PM_7_to_8_2[0] ), .B(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[0] ), .Y(n2489) );
  CLKNAND2X4 U2848 ( .A(n2430), .B(n2414), .Y(n1237) );
  CLKBUFX2 U2853 ( .A(n671), .Y(n3020) );
  BUFX2 U2865 ( .A(n725), .Y(n3021) );
  OAI21X4 U2866 ( .A0(n2211), .A1(n2210), .B0(n2209), .Y(n2224) );
  CLKNAND2X2 U2868 ( .A(n2209), .B(n2219), .Y(n1997) );
  NAND2X3 U2869 ( .A(n2172), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_4[0] ), .Y(
        n1129) );
  INVX1 U2871 ( .A(n2338), .Y(n2334) );
  AND2X4 U2873 ( .A(n2628), .B(n2626), .Y(n995) );
  CLKAND2X2 U2875 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_1[2] ), .B(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[1] ), .Y(n1288) );
  NAND2X5 U2876 ( .A(n2417), .B(n1257), .Y(n1209) );
  NAND2X3 U2881 ( .A(n2272), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[3] ), .Y(
        n2284) );
  CLKNAND2X2 U2884 ( .A(n1195), .B(n2406), .Y(n2366) );
  OAI21X2 U2885 ( .A0(\decoder/u_ACS_matrix/w_PM_5_to_6_3[1] ), .A1(n984), 
        .B0(n2223), .Y(n2308) );
  NAND2BXL U2886 ( .AN(\decoder/w_PM_1[1] ), .B(n671), .Y(n2888) );
  CLKINVX4 U2887 ( .A(n2361), .Y(n957) );
  INVXL U2888 ( .A(n2667), .Y(n3022) );
  INVX2 U2894 ( .A(n2582), .Y(n1279) );
  INVXL U2895 ( .A(n1195), .Y(n3023) );
  CLKNAND2X4 U2899 ( .A(n2646), .B(n1177), .Y(n1246) );
  NAND2BX4 U2900 ( .AN(n2789), .B(n2788), .Y(n2746) );
  CLKINVX2 U2901 ( .A(n2552), .Y(n2553) );
  CLKNAND2X4 U2902 ( .A(n2771), .B(n2791), .Y(n2760) );
  INVX1 U2903 ( .A(n2586), .Y(n1142) );
  NAND3X3 U2904 ( .A(n2628), .B(n2626), .C(n2627), .Y(n2635) );
  OAI22XL U2907 ( .A0(n683), .A1(n2869), .B0(n2834), .B1(n684), .Y(n2825) );
  OAI2B2XL U2908 ( .A1N(\decoder/w_PM_1[3] ), .A0(n683), .B0(n684), .B1(n2892), 
        .Y(n2806) );
  OAI22XL U2909 ( .A0(n684), .A1(n2890), .B0(n2891), .B1(n683), .Y(n2821) );
  INVX3 U2911 ( .A(n2366), .Y(n2367) );
  AOI22X1 U2912 ( .A0(n2909), .A1(n2908), .B0(n2907), .B1(n2906), .Y(n2910) );
  CLKNAND2X12 U2913 ( .A(n1609), .B(n1255), .Y(n2473) );
  INVX8 U2916 ( .A(n1608), .Y(n1609) );
  INVX6 U2918 ( .A(n2473), .Y(n2484) );
  NAND2X3 U2923 ( .A(n2346), .B(n1197), .Y(n1196) );
  MXI2XL U2925 ( .A(n3003), .B(n2641), .S0(n1623), .Y(n735) );
  XOR2X8 U2926 ( .A(n2182), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_3[2] ), .Y(
        n2385) );
  INVXL U2929 ( .A(n2539), .Y(n3026) );
  INVX2 U2931 ( .A(n3026), .Y(n3027) );
  INVX4 U2932 ( .A(n2539), .Y(n2442) );
  INVX3 U2938 ( .A(n2342), .Y(n2412) );
  MXI2XL U2946 ( .A(n2944), .B(n2943), .S0(n2955), .Y(n814) );
  MXI2XL U2947 ( .A(n2299), .B(n2298), .S0(n2955), .Y(n812) );
  MXI2XL U2948 ( .A(n2928), .B(n2927), .S0(n2955), .Y(n813) );
  MXI2XL U2951 ( .A(n2293), .B(n2325), .S0(n2955), .Y(n806) );
  MXI2XL U2952 ( .A(n1009), .B(n2316), .S0(n2955), .Y(n808) );
  MXI2XL U2953 ( .A(n2321), .B(n1232), .S0(n2955), .Y(n810) );
  INVXL U2955 ( .A(n1152), .Y(n3028) );
  INVX2 U2958 ( .A(n3028), .Y(n3029) );
  CLKNAND2X12 U2959 ( .A(n1122), .B(n2178), .Y(n2169) );
  INVXL U2961 ( .A(n2742), .Y(n3030) );
  NAND2X1 U2963 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_1[3] ), .B(
        \decoder/u_ACS_matrix/w_PM_6_to_7_1[4] ), .Y(n1194) );
  CLKNAND2X2 U2964 ( .A(n2608), .B(n2607), .Y(n2618) );
  NOR2X2 U2965 ( .A(n2607), .B(n2362), .Y(n2363) );
  OAI21XL U2966 ( .A0(n2668), .A1(n2721), .B0(n2739), .Y(n2669) );
  CLKAND2X2 U2968 ( .A(n2955), .B(\decoder/u_ACS_matrix/w_data_5_to_6_2[1] ), 
        .Y(n1165) );
  AOI21X6 U2970 ( .A0(n2587), .A1(n1155), .B0(n2586), .Y(n2601) );
  OAI21X4 U2972 ( .A0(n2588), .A1(\decoder/u_ACS_matrix/w_PM_6_to_7_2[4] ), 
        .B0(n2595), .Y(n2642) );
  NOR2X2 U2975 ( .A(n2606), .B(n1095), .Y(n2588) );
  NAND2X3 U2976 ( .A(n2438), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_2[4] ), .Y(
        n2461) );
  OAI21X3 U2979 ( .A0(n2211), .A1(\decoder/u_ACS_matrix/w_PM_5_to_6_2[0] ), 
        .B0(n2257), .Y(n2322) );
  INVX4 U2994 ( .A(\decoder/u_ACS_matrix/w_PM_7_to_8_2[0] ), .Y(n1211) );
  INVX3 U3000 ( .A(n3082), .Y(n2768) );
  INVX1 U3002 ( .A(\decoder/u_ACS_matrix/w_PM_6_to_7_4[1] ), .Y(n1316) );
  CLKMX2X4 U3003 ( .A(n1325), .B(n1323), .S0(n3032), .Y(n1003) );
  MXI2XL U3004 ( .A(n1094), .B(n1097), .S0(n3032), .Y(n3088) );
  OAI22XL U3005 ( .A0(n1098), .A1(n671), .B0(n2824), .B1(n670), .Y(n2819) );
  MXI2X1 U3006 ( .A(n2410), .B(n2409), .S0(n1120), .Y(n762) );
  NOR2BX2 U3007 ( .AN(n1120), .B(n2968), .Y(n769) );
  MXI2XL U3011 ( .A(n2959), .B(n2960), .S0(n1120), .Y(n768) );
  MXI2XL U3012 ( .A(n2406), .B(n3023), .S0(n1120), .Y(n760) );
  MXI2XL U3014 ( .A(n2404), .B(n2403), .S0(n1120), .Y(n759) );
  MXI2XL U3015 ( .A(n2795), .B(n1170), .S0(n1120), .Y(n765) );
  MXI2XL U3016 ( .A(n2948), .B(n1172), .S0(n1120), .Y(n767) );
  MXI2XL U3041 ( .A(n2932), .B(n1171), .S0(n1120), .Y(n766) );
  NAND3X3 U3043 ( .A(n3025), .B(n2255), .C(
        \decoder/u_ACS_matrix/w_PM_5_to_6_1[0] ), .Y(n2252) );
  NAND4X2 U3056 ( .A(n1233), .B(n3034), .C(n2911), .D(n2910), .Y(n2913) );
  OA22X4 U3065 ( .A0(n2883), .A1(\decoder/w_PM_1[6] ), .B0(n2880), .B1(n2879), 
        .Y(n3034) );
  XNOR2X4 U3066 ( .A(n2665), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_4[3] ), .Y(
        n2703) );
  NAND3X4 U3067 ( .A(n973), .B(n988), .C(n3085), .Y(n2665) );
  NOR2X4 U3068 ( .A(n1136), .B(n2321), .Y(n3035) );
  INVX6 U3070 ( .A(n1613), .Y(n1249) );
  NAND2BX1 U3072 ( .AN(\decoder/u_ACS_matrix/w_PM_6_to_7_1[0] ), .B(n2340), 
        .Y(n2343) );
  INVXL U3076 ( .A(n2796), .Y(n3036) );
  INVX1 U3087 ( .A(n3036), .Y(n3037) );
  CLKNAND2X2 U3088 ( .A(n2756), .B(n2757), .Y(n1254) );
  CLKAND2X2 U3090 ( .A(n2597), .B(\decoder/u_ACS_matrix/w_PM_6_to_7_2[0] ), 
        .Y(n1189) );
  AND2X4 U3091 ( .A(n2407), .B(n957), .Y(n2347) );
  MXI2XL U3094 ( .A(n2408), .B(n2407), .S0(n1120), .Y(n761) );
  NAND3X4 U3096 ( .A(n725), .B(n724), .C(n1301), .Y(n1300) );
  BUFX2 U3097 ( .A(n724), .Y(n3066) );
  INVXL U3101 ( .A(io_rst), .Y(n3038) );
  INVX2 U3107 ( .A(n3038), .Y(n3039) );
  CLKBUFX4 U3108 ( .A(n3039), .Y(n1635) );
  NAND2BX4 U3196 ( .AN(n344), .B(n3065), .Y(n2721) );
  MXI2X6 U3197 ( .A(n1569), .B(n1567), .S0(n1565), .Y(n724) );
  OAI2BB1X4 U3199 ( .A0N(n2652), .A1N(n1072), .B0(n1293), .Y(n1127) );
  BUFX12 U3201 ( .A(n2722), .Y(n3067) );
  CLKINVX4 U3202 ( .A(n2714), .Y(n3068) );
  NAND2BX4 U3203 ( .AN(\decoder/u_ACS_matrix/w_PM_7_to_8_3[3] ), .B(n3068), 
        .Y(n2744) );
  BUFX10 U3207 ( .A(n2732), .Y(n3081) );
  INVX2 U3218 ( .A(n3074), .Y(\decoder/w_data_4[4] ) );
  INVX2 U3220 ( .A(n3076), .Y(\decoder/w_data_4[5] ) );
  INVX2 U3223 ( .A(n3078), .Y(\decoder/w_data_4[6] ) );
  AND2X6 U3227 ( .A(n2735), .B(n2723), .Y(n2714) );
  NAND2X2 U3232 ( .A(n2762), .B(n2761), .Y(n3082) );
  OAI21X1 U3233 ( .A0(n2779), .A1(n2744), .B0(n2745), .Y(n1200) );
  NAND3X6 U3234 ( .A(n2778), .B(n2777), .C(n2776), .Y(n2796) );
  NAND2X8 U3235 ( .A(n2796), .B(n2797), .Y(n2981) );
  NAND3X6 U3236 ( .A(n2760), .B(n2748), .C(n3083), .Y(n2797) );
  NOR2BX8 U3237 ( .AN(n2773), .B(n3084), .Y(n3083) );
  INVX4 U3238 ( .A(n1174), .Y(n3084) );
  NAND3X4 U3240 ( .A(n2757), .B(n2756), .C(n1148), .Y(n2763) );
  OAI2BB1X2 U3241 ( .A0N(n2779), .A1N(n2781), .B0(n1200), .Y(n2757) );
  OAI2BB1X1 U3242 ( .A0N(n2982), .A1N(n3086), .B0(n3087), .Y(
        \decoder/u_cmp_sel/N43 ) );
  MXI2X2 U3243 ( .A(n1097), .B(n1094), .S0(n3007), .Y(n3086) );
  MX2X3 U3244 ( .A(n1097), .B(n1094), .S0(n1327), .Y(n2968) );
  CLKINVX16 U3245 ( .A(n1462), .Y(n2938) );
  DFFRQX1 R_160 ( .D(n732), .CK(io_clk), .RN(n1631), .Q(n1436) );
  SNPS_CLOCK_GATE_HIGH_input_fifo_7 \decoder/u_input_shifter/u_input_fifo/clk_gate_data_out_5_reg  ( 
        .CLK(io_clk), .EN(n952), .ENCLK(
        \decoder/u_input_shifter/u_input_fifo/net6035 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_input_fifo_6 \decoder/u_input_shifter/u_input_fifo/clk_gate_data_out_4_reg  ( 
        .CLK(io_clk), .EN(n949), .ENCLK(
        \decoder/u_input_shifter/u_input_fifo/net6030 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_input_fifo_5 \decoder/u_input_shifter/u_input_fifo/clk_gate_data_out_3_reg  ( 
        .CLK(io_clk), .EN(n948), .ENCLK(
        \decoder/u_input_shifter/u_input_fifo/net6025 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_input_fifo_4 \decoder/u_input_shifter/u_input_fifo/clk_gate_data_out_2_reg  ( 
        .CLK(io_clk), .EN(n953), .ENCLK(
        \decoder/u_input_shifter/u_input_fifo/net6020 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_input_fifo_3 \decoder/u_input_shifter/u_input_fifo/clk_gate_data_out_1_reg  ( 
        .CLK(io_clk), .EN(\decoder/u_input_shifter/u_input_fifo/N8 ), .ENCLK(
        \decoder/u_input_shifter/u_input_fifo/net6015 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_input_fifo_2 \decoder/u_input_shifter/u_input_fifo/clk_gate_data_out_8_reg  ( 
        .CLK(io_clk), .EN(\decoder/u_input_shifter/u_input_fifo/N28 ), .ENCLK(
        \decoder/u_input_shifter/u_input_fifo/net6010 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_input_fifo_1 \decoder/u_input_shifter/u_input_fifo/clk_gate_data_out_7_reg  ( 
        .CLK(io_clk), .EN(n950), .ENCLK(
        \decoder/u_input_shifter/u_input_fifo/net6005 ), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_input_fifo_0 \decoder/u_input_shifter/u_input_fifo/clk_gate_data_out_6_reg  ( 
        .CLK(io_clk), .EN(n951), .ENCLK(
        \decoder/u_input_shifter/u_input_fifo/net5999 ), .TE(1'b0) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/PM_out_reg[2]  ( 
        .D(n737), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1627), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[2] ) );
  SDFFRQX4 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/data_out_reg[2]  ( 
        .D(n744), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_data_7_to_8_3[2] ) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_3/u_MEM/PM_out_reg[0]  ( 
        .D(n739), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1628), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_3[0] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/data_out_reg[2]  ( 
        .D(n1165), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_data_6_to_7_1[2] ) );
  SDFFRHQX8 R_254 ( .D(n1112), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), 
        .Q(n2178) );
  SDFFSQX2 R_124 ( .D(n2711), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1482) );
  SDFFRX1 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_4/u_MEM/data_out_reg[1]  ( 
        .D(n1462), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(io_rst), .QN(n1780)
         );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_4/u_MEM/PM_out_reg[6]  ( 
        .D(n720), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(io_rst), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_4[6] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_3/u_MEM/PM_out_reg[1]  ( 
        .D(n935), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1633), .Q(
        \decoder/u_ACS_matrix/w_PM_2_to_3_3[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_3/u_MEM/PM_out_reg[0]  ( 
        .D(n936), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1632), .Q(
        \decoder/u_ACS_matrix/w_PM_2_to_3_3[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_1/u_MEM/PM_out_reg[1]  ( 
        .D(n942), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_2_to_3_1[1] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_4/u_MEM/PM_out_reg[2]  ( 
        .D(n900), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_3_to_4_4[2] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_4/u_MEM/PM_out_reg[0]  ( 
        .D(n932), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1631), .Q(
        \decoder/u_ACS_matrix/w_PM_2_to_3_4[0] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_2/u_MEM/PM_out_reg[4]  ( 
        .D(n839), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1630), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_2[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_5/u_ACS_mem_4/u_MEM/PM_out_reg[4]  ( 
        .D(n818), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_5_to_6_4[4] ) );
  SDFFRHQX2 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_2/u_MEM/PM_out_reg[0]  ( 
        .D(n939), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1626), .Q(
        \decoder/u_ACS_matrix/w_PM_2_to_3_2[0] ) );
  SDFFRX4 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_2/u_MEM/PM_out_reg[5]  ( 
        .D(n794), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(io_rst), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_2[5] ), .QN(n2594) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_7/u_ACS_mem_1/u_MEM/PM_out_reg[6]  ( 
        .D(n1116), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(io_rst), .Q(
        \decoder/u_ACS_matrix/w_PM_7_to_8_1[6] ) );
  SDFFRQX2 \decoder/u_ACS_matrix/u_ACS_col_2/u_ACS_mem_2/u_MEM/PM_out_reg[1]  ( 
        .D(n938), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1634), .Q(
        \decoder/u_ACS_matrix/w_PM_2_to_3_2[1] ) );
  SDFFRHQX4 \decoder/u_ACS_matrix/u_ACS_col_3/u_ACS_mem_4/u_MEM/data_out_reg[2]  ( 
        .D(n903), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(io_rst), .Q(
        \decoder/u_ACS_matrix/w_data_3_to_4_4[2] ) );
  SDFFSX2 R_224 ( .D(n1869), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(io_rst), 
        .Q(n1349) );
  SDFFRQX2 R_203 ( .D(n2522), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(io_rst), 
        .Q(n1381) );
  SDFFSX1 R_285 ( .D(n2938), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(io_rst), 
        .Q(n1097), .QN(n732) );
  SDFFSHQX2 R_57 ( .D(n2789), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1544) );
  SDFFSHQX1 R_102 ( .D(n2306), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1633), 
        .Q(n1502) );
  SDFFSHQX4 R_103 ( .D(n2305), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1629), 
        .Q(n1500) );
  SDFFRHQX8 \decoder/u_ACS_matrix/u_ACS_col_6/u_ACS_mem_1/u_MEM/PM_out_reg[4]  ( 
        .D(n807), .SI(1'b0), .SE(1'b0), .CK(io_clk), .RN(n1629), .Q(
        \decoder/u_ACS_matrix/w_PM_6_to_7_1[4] ) );
  SDFFSHQX1 R_71 ( .D(n1132), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1530) );
  SDFFSHQX4 R_67 ( .D(n2781), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1626), 
        .Q(n1536) );
  SDFFSHQX2 R_236 ( .D(n2698), .SI(1'b0), .SE(1'b0), .CK(io_clk), .SN(n1635), 
        .Q(n1336) );
  BUFX14 U1101 ( .A(n2965), .Y(n1120) );
  CLKNAND2X2 U1104 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_3[0] ), .B(n1804), 
        .Y(n1863) );
  INVX2 U1128 ( .A(n2151), .Y(n2123) );
  BUFX2 U1134 ( .A(n2151), .Y(n3069) );
  OAI21X8 U1146 ( .A0(n2130), .A1(n2129), .B0(n2128), .Y(n2954) );
  MX2X2 U1161 ( .A(n2118), .B(n2166), .S0(n2128), .Y(n783) );
  CLKNAND2X8 U1176 ( .A(n2126), .B(n2150), .Y(n2128) );
  OAI21X6 U1189 ( .A0(n2130), .A1(n2129), .B0(n2128), .Y(n3089) );
  AOI21X6 U1191 ( .A0(n2114), .A1(n2115), .B0(n2113), .Y(n2130) );
  CLKAND2X2 U1213 ( .A(n3089), .B(\decoder/u_ACS_matrix/w_data_5_to_6_2[1] ), 
        .Y(n792) );
  NOR2X1 U1231 ( .A(n2703), .B(n2682), .Y(n1037) );
  AOI21X2 U1232 ( .A0(n2682), .A1(n2703), .B0(n2704), .Y(n2674) );
  NAND3X3 U1238 ( .A(n1318), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[1] ), .C(
        n1317), .Y(n2678) );
  XNOR2X2 U1247 ( .A(n1048), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[5] ), .Y(
        n2700) );
  INVX3 U1250 ( .A(n2312), .Y(n1160) );
  NAND2X6 U1252 ( .A(n1161), .B(n2292), .Y(n1287) );
  INVX1 U1258 ( .A(n2284), .Y(n1290) );
  OAI21XL U1260 ( .A0(n2676), .A1(\decoder/u_ACS_matrix/w_PM_7_to_8_3[3] ), 
        .B0(n2673), .Y(n2704) );
  NOR2X3 U1264 ( .A(n2678), .B(n1202), .Y(n2676) );
  NOR2X4 U1300 ( .A(n2688), .B(n2702), .Y(n2691) );
  OAI21X4 U1305 ( .A0(n2211), .A1(n2210), .B0(n2225), .Y(n1999) );
  OAI2B1XL U1338 ( .A1N(n1620), .A0(n2160), .B0(n1064), .Y(n772) );
  OAI2B1XL U1339 ( .A1N(n2161), .A0(n2163), .B0(n2162), .Y(n1064) );
  NAND2X4 U1353 ( .A(n2160), .B(n2162), .Y(n2163) );
  NOR2X3 U1387 ( .A(n1992), .B(n1274), .Y(n1993) );
  AOI21X4 U1416 ( .A0(n2146), .A1(n2145), .B0(n1995), .Y(n2006) );
  NAND2X2 U1421 ( .A(n1613), .B(n1248), .Y(n2209) );
  NAND2X2 U1425 ( .A(n2675), .B(n2674), .Y(n2687) );
  NAND2X8 U1446 ( .A(n2663), .B(n2660), .Y(n2679) );
  NAND2X3 U1511 ( .A(n2661), .B(n2679), .Y(n2698) );
  INVX1 U1513 ( .A(n2225), .Y(n2228) );
  NOR2BX8 U1515 ( .AN(n2222), .B(n2220), .Y(n2221) );
  AOI2BB1X2 U1521 ( .A0N(n2222), .A1N(\decoder/u_ACS_matrix/w_PM_5_to_6_4[1] ), 
        .B0(n2221), .Y(n2307) );
  OAI21BX4 U1553 ( .A0(n2665), .A1(n1219), .B0N(
        \decoder/u_ACS_matrix/w_PM_7_to_8_4[4] ), .Y(n2661) );
  AND2X4 U1594 ( .A(n2681), .B(n2680), .Y(n2672) );
  AOI21X3 U1603 ( .A0(n2300), .A1(n2214), .B0(n2326), .Y(n2239) );
  NOR2X4 U1612 ( .A(n2328), .B(n2327), .Y(n2326) );
  MXI2X2 U1623 ( .A(n2311), .B(n2310), .S0(n2964), .Y(n799) );
  INVX1 U1624 ( .A(n2274), .Y(n2319) );
  NAND2X4 U1625 ( .A(n2345), .B(n1193), .Y(n2349) );
  CLKINVX2 U1666 ( .A(n2765), .Y(n2784) );
  NAND3X2 U1674 ( .A(n1228), .B(n2598), .C(n998), .Y(n2600) );
  CLKNAND2X2 U1687 ( .A(n1228), .B(n2343), .Y(n2650) );
  INVXL U1721 ( .A(n2738), .Y(n2668) );
  CLKNAND2X2 U1723 ( .A(n2666), .B(n2786), .Y(n2738) );
  NOR2X6 U1728 ( .A(n2716), .B(n2715), .Y(n2772) );
  MXI2X4 U1772 ( .A(n2734), .B(n1205), .S0(n2733), .Y(n2741) );
  XNOR2X4 U1784 ( .A(n2506), .B(n2505), .Y(n2511) );
  CLKINVX3 U1818 ( .A(n2477), .Y(n2506) );
  INVX4 U1848 ( .A(n2714), .Y(n2716) );
  CLKINVX2 U1852 ( .A(n2749), .Y(n2750) );
  CLKNAND2X2 U1906 ( .A(n2746), .B(n2747), .Y(n2756) );
  BUFX8 U1925 ( .A(n2769), .Y(n1148) );
  OR2X1 U1938 ( .A(n725), .B(n724), .Y(n2728) );
  INVX2 U1947 ( .A(n2781), .Y(n2743) );
  NOR2X4 U1952 ( .A(n3006), .B(n2321), .Y(n2275) );
  CLKNAND2X2 U1956 ( .A(n1795), .B(n1794), .Y(n1776) );
  NOR2BXL U1959 ( .AN(\decoder/u_ACS_matrix/w_data_3_to_4_2[1] ), .B(n1132), 
        .Y(n876) );
  OAI2B2X2 U1970 ( .A1N(n1743), .A0(n1735), .B0(n1734), .B1(n1746), .Y(n1750)
         );
  CLKINVX2 U1973 ( .A(n1743), .Y(n1836) );
  AOI2BB2X4 U1985 ( .B0(n1745), .B1(n1744), .A0N(n1743), .A1N(n1835), .Y(n1749) );
  OAI2BB1X4 U1996 ( .A0N(n1868), .A1N(n3090), .B0(n1869), .Y(n1876) );
  CLKINVX40 U2015 ( .A(\decoder/u_ACS_matrix/w_PM_3_to_4_3[2] ), .Y(n3090) );
  INVX1 U2027 ( .A(n1881), .Y(n1885) );
  INVX6 U2038 ( .A(n1834), .Y(n2936) );
  OAI21X3 U2099 ( .A0(n891), .A1(n986), .B0(n2019), .Y(n2082) );
  AOI22X1 U2114 ( .A0(n1926), .A1(n1928), .B0(n1874), .B1(n1930), .Y(n1878) );
  NAND2X3 U2127 ( .A(n2043), .B(n2042), .Y(n2046) );
  AOI2BB2X1 U2128 ( .B0(n1922), .B1(n1876), .A0N(n1879), .A1N(n1880), .Y(n1877) );
  MXI2X1 U2173 ( .A(n1963), .B(n1962), .S0(n1958), .Y(n831) );
  NAND2BX4 U2191 ( .AN(n1962), .B(n1963), .Y(n1852) );
  NOR2X1 U2226 ( .A(n1804), .B(n1799), .Y(n3091) );
  NOR2X2 U2255 ( .A(n1804), .B(n1799), .Y(n1898) );
  NOR2X6 U2266 ( .A(n2103), .B(n2100), .Y(n3012) );
  OAI2BB1X4 U2323 ( .A0N(n2103), .A1N(n2100), .B0(n963), .Y(n2148) );
  INVX3 U2330 ( .A(\decoder/u_ACS_matrix/w_PM_5_to_6_2[2] ), .Y(n2100) );
  AOI21X6 U2387 ( .A0(n2157), .A1(n2159), .B0(n2104), .Y(n2115) );
  OAI2BB1X2 U2408 ( .A0N(n2166), .A1N(n2121), .B0(n2152), .Y(n2126) );
  OAI21X1 U2418 ( .A0(n2154), .A1(n2152), .B0(n3069), .Y(n2155) );
  NAND2X2 U2421 ( .A(n2125), .B(n2151), .Y(n2152) );
  NAND2X6 U2436 ( .A(n2150), .B(n2124), .Y(n2129) );
  OAI2BB1X2 U2445 ( .A0N(n2688), .A1N(n2702), .B0(n2696), .Y(n1292) );
  BUFX2 U2454 ( .A(n749), .Y(n2989) );
  CLKINVX3 U2455 ( .A(n749), .Y(n2414) );
  AOI2BB1X1 U2465 ( .A0N(n2226), .A1N(n2209), .B0(n1996), .Y(n2003) );
  NAND2X2 U2489 ( .A(n2233), .B(n2305), .Y(n2234) );
  OAI2BB1X4 U2493 ( .A0N(n2218), .A1N(n2223), .B0(n2217), .Y(n2305) );
  XNOR2X4 U2524 ( .A(n973), .B(n2734), .Y(n2670) );
  AOI21X1 U2613 ( .A0(n2708), .A1(n2670), .B0(n2669), .Y(n2683) );
  NOR2X1 U2626 ( .A(n2250), .B(\decoder/u_ACS_matrix/w_PM_5_to_6_1[1] ), .Y(
        n2253) );
  NAND3X2 U2644 ( .A(n2695), .B(n2694), .C(n2693), .Y(n2696) );
  NOR2X8 U2697 ( .A(n2658), .B(n2659), .Y(n2660) );
  NAND2X4 U2722 ( .A(n3021), .B(n3066), .Y(n2658) );
  BUFX14 U2724 ( .A(n2969), .Y(n1623) );
  NAND2BX8 U2735 ( .AN(n2724), .B(n3081), .Y(n2663) );
  INVX3 U2738 ( .A(n2641), .Y(n2622) );
  CLKNAND2X2 U2743 ( .A(n1208), .B(n2481), .Y(n2477) );
  NAND2X4 U2744 ( .A(n1126), .B(n1004), .Y(n3092) );
  NAND2X4 U2836 ( .A(n1126), .B(n1004), .Y(n2977) );
  BUFX2 U2867 ( .A(n725), .Y(n3085) );
  BUFX5 U2880 ( .A(n725), .Y(n1205) );
  MXI2X1 U2891 ( .A(n2651), .B(n2650), .S0(n1623), .Y(n739) );
  MXI2XL U2893 ( .A(n1172), .B(n2948), .S0(n1623), .Y(n742) );
  MXI2XL U2896 ( .A(n1170), .B(n2795), .S0(n1623), .Y(n740) );
  MXI2XL U2897 ( .A(n2960), .B(n2959), .S0(n1623), .Y(n743) );
  MXI2XL U2898 ( .A(n1171), .B(n2932), .S0(n1623), .Y(n741) );
  MXI2XL U2905 ( .A(n2644), .B(n2643), .S0(n1623), .Y(n736) );
  INVXL U2928 ( .A(n2648), .Y(n3093) );
  INVX2 U2930 ( .A(n3093), .Y(n3094) );
  INVX3 U2936 ( .A(n2779), .Y(n2742) );
  CLKNAND2X4 U2943 ( .A(n2783), .B(n2765), .Y(n2773) );
  XOR2X8 U2962 ( .A(n2753), .B(\decoder/u_ACS_matrix/w_PM_7_to_8_3[6] ), .Y(
        n2783) );
  AOI21X6 U2971 ( .A0(n2775), .A1(n2785), .B0(n2774), .Y(n2776) );
  AOI21X1 U2978 ( .A0(n2754), .A1(n1148), .B0(n2790), .Y(n3095) );
  NAND2X2 U2981 ( .A(n2202), .B(n2384), .Y(n1063) );
  CLKNAND2X4 U2982 ( .A(n1263), .B(n1262), .Y(n2197) );
  NAND2X5 U2985 ( .A(n2173), .B(n994), .Y(n2386) );
  AOI21X2 U3001 ( .A0(n2754), .A1(n1148), .B0(n2790), .Y(n2761) );
  CLKINVX6 U3019 ( .A(n2656), .Y(n2592) );
  CLKNAND2X4 U3020 ( .A(n2613), .B(n2656), .Y(n2627) );
  MXI2XL U3021 ( .A(n2657), .B(n2656), .S0(n1623), .Y(n734) );
  NAND2X4 U3022 ( .A(n1256), .B(n2473), .Y(n2417) );
  OAI21X1 U3042 ( .A0(n2648), .A1(n2647), .B0(n1246), .Y(n3096) );
  OAI21X4 U3069 ( .A0(n2648), .A1(n2647), .B0(n1246), .Y(n2617) );
  CLKNAND2X4 U3071 ( .A(n2413), .B(n2650), .Y(n2614) );
  NOR2X4 U3073 ( .A(n2341), .B(n2413), .Y(n2605) );
  INVXL U3075 ( .A(n2413), .Y(n2651) );
  OAI2B1X2 U3095 ( .A1N(n2731), .A0(\decoder/u_ACS_matrix/w_PM_7_to_8_4[4] ), 
        .B0(n2749), .Y(n2790) );
  NAND3X3 U3100 ( .A(n1218), .B(n1217), .C(
        \decoder/u_ACS_matrix/w_PM_7_to_8_4[3] ), .Y(n2731) );
  AND2X4 U3103 ( .A(n1015), .B(n1016), .Y(n2759) );
  NAND2X2 U3112 ( .A(n2743), .B(n2742), .Y(n1015) );
  CLKNAND2X8 U3113 ( .A(n2523), .B(n2522), .Y(n2710) );
  NAND3BX2 U3114 ( .AN(n724), .B(n2732), .C(n2737), .Y(n2730) );
  INVX2 U3115 ( .A(n2786), .Y(n2667) );
  INVXL U3165 ( .A(n2579), .Y(n3097) );
  INVX2 U3168 ( .A(n3097), .Y(n3098) );
  BUFX3 U3208 ( .A(n2340), .Y(n1198) );
endmodule

