module ACS_matrix(clk,
				  rst,
				  data_id,
				  input_valid,
				  data_recv_1,
				  data_recv_2,
				  data_recv_3,
				  data_recv_4,
				  data_recv_5,
				  data_recv_6,
				  data_recv_7,
				  data_recv_8,
				  bus_sig_1,
				  bus_sig_2,
				  bus_sig_3,
				  bus_sig_4,
				  bus_sig_5,
				  bus_sig_6,
				  bus_sig_7,
				  bus_sig_8,
				  PM_8_1,
				  PM_8_2,
				  PM_8_3,
				  PM_8_4);
	
	input clk,rst,input_valid;
	input [1:0] data_recv_1,data_recv_2,data_recv_3,data_recv_4,data_recv_5,data_recv_6,data_recv_7,data_recv_8;
	input [2:0] data_id;

	output [6:0] PM_8_1,PM_8_2,PM_8_3,PM_8_4;
	output [14:0] bus_sig_1,bus_sig_2,bus_sig_3,bus_sig_4,bus_sig_5,bus_sig_6,bus_sig_7,bus_sig_8;

	//reg [1:0] addr_init_1,addr_init_2,addr_init_3,addr_init_4;
	//reg [6:0] PM_init;

	wire dec_out_1_1,dec_out_1_2,dec_out_1_3,dec_out_1_4,
		 dec_out_2_1,dec_out_2_2,dec_out_2_3,dec_out_2_4,
		 dec_out_3_1,dec_out_3_2,dec_out_3_3,dec_out_3_4,
		 dec_out_4_1,dec_out_4_2,dec_out_4_3,dec_out_4_4,
		 dec_out_5_1,dec_out_5_2,dec_out_5_3,dec_out_5_4,
		 dec_out_6_1,dec_out_6_2,dec_out_6_3,dec_out_6_4,
		 dec_out_7_1,dec_out_7_2,dec_out_7_3,dec_out_7_4,
		 dec_out_8_1,dec_out_8_2,dec_out_8_3,dec_out_8_4,
		 data_rdy;

	wire [1:0] addr_1_to_2_1,addr_1_to_2_2,addr_1_to_2_3,addr_1_to_2_4,
			   addr_2_to_3_1,addr_2_to_3_2,addr_2_to_3_3,addr_2_to_3_4,
			   addr_3_to_4_1,addr_3_to_4_2,addr_3_to_4_3,addr_3_to_4_4,
			   addr_4_to_5_1,addr_4_to_5_2,addr_4_to_5_3,addr_4_to_5_4,
			   addr_5_to_6_1,addr_5_to_6_2,addr_5_to_6_3,addr_5_to_6_4,
			   addr_6_to_7_1,addr_6_to_7_2,addr_6_to_7_3,addr_6_to_7_4,
			   addr_7_to_8_1,addr_7_to_8_2,addr_7_to_8_3,addr_7_to_8_4,
			   w_addr_8_1,w_addr_8_2,w_addr_8_3,w_addr_8_4;

	wire [2:0] data_id_1_to_2,data_id_2_to_3,data_id_3_to_4,data_id_4_to_5,data_id_5_to_6,data_id_6_to_7,data_id_7_to_8,w_data_id_8;

	wire [6:0] PM_1_to_2_1,PM_1_to_2_2,PM_1_to_2_3,PM_1_to_2_4,
			   PM_2_to_3_1,PM_2_to_3_2,PM_2_to_3_3,PM_2_to_3_4,
			   PM_3_to_4_1,PM_3_to_4_2,PM_3_to_4_3,PM_3_to_4_4,
			   PM_4_to_5_1,PM_4_to_5_2,PM_4_to_5_3,PM_4_to_5_4,
			   PM_5_to_6_1,PM_5_to_6_2,PM_5_to_6_3,PM_5_to_6_4,
			   PM_6_to_7_1,PM_6_to_7_2,PM_6_to_7_3,PM_6_to_7_4,
			   PM_7_to_8_1,PM_7_to_8_2,PM_7_to_8_3,PM_7_to_8_4;


	//always begin
	//	addr_init_1 = 2'b00;
	//	addr_init_2 = 2'b01;
	//	addr_init_3 = 2'b10;
	//	addr_init_4 = 2'b11;
	//	PM_init = 7'b0000000;
	//end

	ACS_col u_ACS_col_1(.clk(clk),
			   .rst(rst),
			   .data_id(data_id),
			   .input_valid(input_valid),
			   .data_recv(data_recv_1),
			   .PM_in_1_1(7'b0000000),
			   .PM_in_1_2(7'b0000000),
			   .PM_in_2_1(7'b0000000),
			   .PM_in_2_2(7'b0000000),
			   .PM_in_3_1(7'b0000000),
			   .PM_in_3_2(7'b0000000),
			   .PM_in_4_1(7'b0000000),
			   .PM_in_4_2(7'b0000000),
			   .addr_in_1_1(2'b00),
			   .addr_in_1_2(2'b00),
			   .addr_in_2_1(2'b01),
			   .addr_in_2_2(2'b01),
			   .addr_in_3_1(2'b10),
			   .addr_in_3_2(2'b10),
			   .addr_in_4_1(2'b11),
			   .addr_in_4_2(2'b11),
			   .addr_out_1(addr_1_to_2_1),
			   .addr_out_2(addr_1_to_2_2),
			   .addr_out_3(addr_1_to_2_3),
			   .addr_out_4(addr_1_to_2_4),
			   .PM_out_1(PM_1_to_2_1),
			   .PM_out_2(PM_1_to_2_2),
			   .PM_out_3(PM_1_to_2_3),
			   .PM_out_4(PM_1_to_2_4),
			   .dec_out_1(dec_out_1_1),
			   .dec_out_2(dec_out_1_2),
			   .dec_out_3(dec_out_1_3),
			   .dec_out_4(dec_out_1_4),
			   .data_id_out(data_id_1_to_2),
			   .data_rdy(data_rdy));

	ACS_col u_ACS_col_2(.clk(clk),
			   .rst(rst),
			   .data_id(data_id_1_to_2),
			   .input_valid(input_valid),
			   .data_recv(data_recv_2),
			   .PM_in_1_1(PM_1_to_2_1),
			   .PM_in_1_2(PM_1_to_2_2),
			   .PM_in_2_1(PM_1_to_2_3),
			   .PM_in_2_2(PM_1_to_2_4),
			   .PM_in_3_1(PM_1_to_2_1),
			   .PM_in_3_2(PM_1_to_2_2),
			   .PM_in_4_1(PM_1_to_2_3),
			   .PM_in_4_2(PM_1_to_2_4),
			   .addr_in_1_1(addr_1_to_2_1),
			   .addr_in_1_2(addr_1_to_2_2),
			   .addr_in_2_1(addr_1_to_2_3),
			   .addr_in_2_2(addr_1_to_2_4),
			   .addr_in_3_1(addr_1_to_2_1),
			   .addr_in_3_2(addr_1_to_2_2),
			   .addr_in_4_1(addr_1_to_2_3),
			   .addr_in_4_2(addr_1_to_2_4),
			   .addr_out_1(addr_2_to_3_1),
			   .addr_out_2(addr_2_to_3_2),
			   .addr_out_3(addr_2_to_3_3),
			   .addr_out_4(addr_2_to_3_4),
			   .PM_out_1(PM_2_to_3_1),
			   .PM_out_2(PM_2_to_3_2),
			   .PM_out_3(PM_2_to_3_3),
			   .PM_out_4(PM_2_to_3_4),
			   .dec_out_1(dec_out_2_1),
			   .dec_out_2(dec_out_2_2),
			   .dec_out_3(dec_out_2_3),
			   .dec_out_4(dec_out_2_4),
			   .data_id_out(data_id_2_to_3),
			   .data_rdy(data_rdy));

	ACS_col u_ACS_col_3(.clk(clk),
			   .rst(rst),
			   .data_id(data_id_2_to_3),
			   .input_valid(input_valid),
			   .data_recv(data_recv_3),
			   .PM_in_1_1(PM_2_to_3_1),
			   .PM_in_1_2(PM_2_to_3_2),
			   .PM_in_2_1(PM_2_to_3_3),
			   .PM_in_2_2(PM_2_to_3_4),
			   .PM_in_3_1(PM_2_to_3_1),
			   .PM_in_3_2(PM_2_to_3_2),
			   .PM_in_4_1(PM_2_to_3_3),
			   .PM_in_4_2(PM_2_to_3_4),
			   .addr_in_1_1(addr_2_to_3_1),
			   .addr_in_1_2(addr_2_to_3_2),
			   .addr_in_2_1(addr_2_to_3_3),
			   .addr_in_2_2(addr_2_to_3_4),
			   .addr_in_3_1(addr_2_to_3_1),
			   .addr_in_3_2(addr_2_to_3_2),
			   .addr_in_4_1(addr_2_to_3_3),
			   .addr_in_4_2(addr_2_to_3_4),
			   .addr_out_1(addr_3_to_4_1),
			   .addr_out_2(addr_3_to_4_2),
			   .addr_out_3(addr_3_to_4_3),
			   .addr_out_4(addr_3_to_4_4),
			   .PM_out_1(PM_3_to_4_1),
			   .PM_out_2(PM_3_to_4_2),
			   .PM_out_3(PM_3_to_4_3),
			   .PM_out_4(PM_3_to_4_4),
			   .dec_out_1(dec_out_3_1),
			   .dec_out_2(dec_out_3_2),
			   .dec_out_3(dec_out_3_3),
			   .dec_out_4(dec_out_3_4),
			   .data_id_out(data_id_3_to_4),
			   .data_rdy(data_rdy));

	ACS_col u_ACS_col_4(.clk(clk),
			   .rst(rst),
			   .data_id(data_id_3_to_4),
			   .input_valid(input_valid),
			   .data_recv(data_recv_4),
			   .PM_in_1_1(PM_3_to_4_1),
			   .PM_in_1_2(PM_3_to_4_2),
			   .PM_in_2_1(PM_3_to_4_3),
			   .PM_in_2_2(PM_3_to_4_4),
			   .PM_in_3_1(PM_3_to_4_1),
			   .PM_in_3_2(PM_3_to_4_2),
			   .PM_in_4_1(PM_3_to_4_3),
			   .PM_in_4_2(PM_3_to_4_4),
			   .addr_in_1_1(addr_3_to_4_1),
			   .addr_in_1_2(addr_3_to_4_2),
			   .addr_in_2_1(addr_3_to_4_3),
			   .addr_in_2_2(addr_3_to_4_4),
			   .addr_in_3_1(addr_3_to_4_1),
			   .addr_in_3_2(addr_3_to_4_2),
			   .addr_in_4_1(addr_3_to_4_3),
			   .addr_in_4_2(addr_3_to_4_4),
			   .addr_out_1(addr_4_to_5_1),
			   .addr_out_2(addr_4_to_5_2),
			   .addr_out_3(addr_4_to_5_3),
			   .addr_out_4(addr_4_to_5_4),
			   .PM_out_1(PM_4_to_5_1),
			   .PM_out_2(PM_4_to_5_2),
			   .PM_out_3(PM_4_to_5_3),
			   .PM_out_4(PM_4_to_5_4),
			   .dec_out_1(dec_out_4_1),
			   .dec_out_2(dec_out_4_2),
			   .dec_out_3(dec_out_4_3),
			   .dec_out_4(dec_out_4_4),
			   .data_id_out(data_id_4_to_5),
			   .data_rdy(data_rdy));

	ACS_col u_ACS_col_5(.clk(clk),
			   .rst(rst),
			   .data_id(data_id_4_to_5),
			   .input_valid(input_valid),
			   .data_recv(data_recv_5),
			   .PM_in_1_1(PM_4_to_5_1),
			   .PM_in_1_2(PM_4_to_5_2),
			   .PM_in_2_1(PM_4_to_5_3),
			   .PM_in_2_2(PM_4_to_5_4),
			   .PM_in_3_1(PM_4_to_5_1),
			   .PM_in_3_2(PM_4_to_5_2),
			   .PM_in_4_1(PM_4_to_5_3),
			   .PM_in_4_2(PM_4_to_5_4),
			   .addr_in_1_1(addr_4_to_5_1),
			   .addr_in_1_2(addr_4_to_5_2),
			   .addr_in_2_1(addr_4_to_5_3),
			   .addr_in_2_2(addr_4_to_5_4),
			   .addr_in_3_1(addr_4_to_5_1),
			   .addr_in_3_2(addr_4_to_5_2),
			   .addr_in_4_1(addr_4_to_5_3),
			   .addr_in_4_2(addr_4_to_5_4),
			   .addr_out_1(addr_5_to_6_1),
			   .addr_out_2(addr_5_to_6_2),
			   .addr_out_3(addr_5_to_6_3),
			   .addr_out_4(addr_5_to_6_4),
			   .PM_out_1(PM_5_to_6_1),
			   .PM_out_2(PM_5_to_6_2),
			   .PM_out_3(PM_5_to_6_3),
			   .PM_out_4(PM_5_to_6_4),
			   .dec_out_1(dec_out_5_1),
			   .dec_out_2(dec_out_5_2),
			   .dec_out_3(dec_out_5_3),
			   .dec_out_4(dec_out_5_4),
			   .data_id_out(data_id_5_to_6),
			   .data_rdy(data_rdy));

	ACS_col u_ACS_col_6(.clk(clk),
			   .rst(rst),
			   .data_id(data_id_5_to_6),
			   .input_valid(input_valid),
			   .data_recv(data_recv_6),
			   .PM_in_1_1(PM_5_to_6_1),
			   .PM_in_1_2(PM_5_to_6_2),
			   .PM_in_2_1(PM_5_to_6_3),
			   .PM_in_2_2(PM_5_to_6_4),
			   .PM_in_3_1(PM_5_to_6_1),
			   .PM_in_3_2(PM_5_to_6_2),
			   .PM_in_4_1(PM_5_to_6_3),
			   .PM_in_4_2(PM_5_to_6_4),
			   .addr_in_1_1(addr_5_to_6_1),
			   .addr_in_1_2(addr_5_to_6_2),
			   .addr_in_2_1(addr_5_to_6_3),
			   .addr_in_2_2(addr_5_to_6_4),
			   .addr_in_3_1(addr_5_to_6_1),
			   .addr_in_3_2(addr_5_to_6_2),
			   .addr_in_4_1(addr_5_to_6_3),
			   .addr_in_4_2(addr_5_to_6_4),
			   .addr_out_1(addr_6_to_7_1),
			   .addr_out_2(addr_6_to_7_2),
			   .addr_out_3(addr_6_to_7_3),
			   .addr_out_4(addr_6_to_7_4),
			   .PM_out_1(PM_6_to_7_1),
			   .PM_out_2(PM_6_to_7_2),
			   .PM_out_3(PM_6_to_7_3),
			   .PM_out_4(PM_6_to_7_4),
			   .dec_out_1(dec_out_6_1),
			   .dec_out_2(dec_out_6_2),
			   .dec_out_3(dec_out_6_3),
			   .dec_out_4(dec_out_6_4),
			   .data_id_out(data_id_6_to_7),
			   .data_rdy(data_rdy));

	ACS_col u_ACS_col_7(.clk(clk),
			   .rst(rst),
			   .data_id(data_id_6_to_7),
			   .input_valid(input_valid),
			   .data_recv(data_recv_7),
			   .PM_in_1_1(PM_6_to_7_1),
			   .PM_in_1_2(PM_6_to_7_2),
			   .PM_in_2_1(PM_6_to_7_3),
			   .PM_in_2_2(PM_6_to_7_4),
			   .PM_in_3_1(PM_6_to_7_1),
			   .PM_in_3_2(PM_6_to_7_2),
			   .PM_in_4_1(PM_6_to_7_3),
			   .PM_in_4_2(PM_6_to_7_4),
			   .addr_in_1_1(addr_6_to_7_1),
			   .addr_in_1_2(addr_6_to_7_2),
			   .addr_in_2_1(addr_6_to_7_3),
			   .addr_in_2_2(addr_6_to_7_4),
			   .addr_in_3_1(addr_6_to_7_1),
			   .addr_in_3_2(addr_6_to_7_2),
			   .addr_in_4_1(addr_6_to_7_3),
			   .addr_in_4_2(addr_6_to_7_4),
			   .addr_out_1(addr_7_to_8_1),
			   .addr_out_2(addr_7_to_8_2),
			   .addr_out_3(addr_7_to_8_3),
			   .addr_out_4(addr_7_to_8_4),
			   .PM_out_1(PM_7_to_8_1),
			   .PM_out_2(PM_7_to_8_2),
			   .PM_out_3(PM_7_to_8_3),
			   .PM_out_4(PM_7_to_8_4),
			   .dec_out_1(dec_out_7_1),
			   .dec_out_2(dec_out_7_2),
			   .dec_out_3(dec_out_7_3),
			   .dec_out_4(dec_out_7_4),
			   .data_id_out(data_id_7_to_8),
			   .data_rdy(data_rdy));

	ACS_col u_ACS_col_8(.clk(clk),
			   .rst(rst),
			   .data_id(data_id_7_to_8),
			   .input_valid(input_valid),
			   .data_recv(data_recv_8),
			   .PM_in_1_1(PM_7_to_8_1),
			   .PM_in_1_2(PM_7_to_8_2),
			   .PM_in_2_1(PM_7_to_8_3),
			   .PM_in_2_2(PM_7_to_8_4),
			   .PM_in_3_1(PM_7_to_8_1),
			   .PM_in_3_2(PM_7_to_8_2),
			   .PM_in_4_1(PM_7_to_8_3),
			   .PM_in_4_2(PM_7_to_8_4),
			   .addr_in_1_1(addr_7_to_8_1),
			   .addr_in_1_2(addr_7_to_8_2),
			   .addr_in_2_1(addr_7_to_8_3),
			   .addr_in_2_2(addr_7_to_8_4),
			   .addr_in_3_1(addr_7_to_8_1),
			   .addr_in_3_2(addr_7_to_8_2),
			   .addr_in_4_1(addr_7_to_8_3),
			   .addr_in_4_2(addr_7_to_8_4),
			   .addr_out_1(w_addr_8_1),
			   .addr_out_2(w_addr_8_2),
			   .addr_out_3(w_addr_8_3),
			   .addr_out_4(w_addr_8_4),
			   .PM_out_1(PM_8_1),
			   .PM_out_2(PM_8_2),
			   .PM_out_3(PM_8_3),
			   .PM_out_4(PM_8_4),
			   .dec_out_1(dec_out_8_1),
			   .dec_out_2(dec_out_8_2),
			   .dec_out_3(dec_out_8_3),
			   .dec_out_4(dec_out_8_4),
			   .data_id_out(w_data_id_8),
			   .data_rdy(data_rdy));

	// assign bus_sig_n = {data_id_n_to_n+1,
	//					   addr_n_to_n+1_4,dec_out_n_4,
	//					   addr_n_to_n+1_3,dec_out_n_3,
	//					   addr_n_to_n+1_2,dec_out_n_2,
	//					   addr_n_to_n+1_1,dec_out_n_1};

	assign bus_sig_1 = {data_id_1_to_2,
						addr_1_to_2_4,dec_out_1_4,
						addr_1_to_2_3,dec_out_1_3,
						addr_1_to_2_2,dec_out_1_2,
						addr_1_to_2_1,dec_out_1_1};
	assign bus_sig_2 = {data_id_2_to_3,
						addr_2_to_3_4,dec_out_2_4,
						addr_2_to_3_3,dec_out_2_3,
						addr_2_to_3_2,dec_out_2_2,
						addr_2_to_3_1,dec_out_2_1};
	assign bus_sig_3 = {data_id_3_to_4,
						addr_3_to_4_4,dec_out_3_4,
						addr_3_to_4_3,dec_out_3_3,
						addr_3_to_4_2,dec_out_3_2,
						addr_3_to_4_1,dec_out_3_1};
	assign bus_sig_4 = {data_id_4_to_5,
						addr_4_to_5_4,dec_out_4_4,
						addr_4_to_5_3,dec_out_4_3,
						addr_4_to_5_2,dec_out_4_2,
						addr_4_to_5_1,dec_out_4_1};
	assign bus_sig_5 = {data_id_5_to_6,
						addr_5_to_6_4,dec_out_5_4,
						addr_5_to_6_3,dec_out_5_3,
						addr_5_to_6_2,dec_out_5_2,
						addr_5_to_6_1,dec_out_5_1};
	assign bus_sig_6 = {data_id_6_to_7,
						addr_6_to_7_4,dec_out_6_4,
						addr_6_to_7_3,dec_out_6_3,
						addr_6_to_7_2,dec_out_6_2,
						addr_6_to_7_1,dec_out_6_1};
	assign bus_sig_7 = {data_id_7_to_8,
						addr_7_to_8_4,dec_out_7_4,
						addr_7_to_8_3,dec_out_7_3,
						addr_7_to_8_2,dec_out_7_2,
						addr_7_to_8_1,dec_out_7_1};
	assign bus_sig_8 = {w_data_id_8,
						w_addr_8_4,dec_out_8_4,
						w_addr_8_3,dec_out_8_3,
						w_addr_8_2,dec_out_8_2,
						w_addr_8_1,dec_out_8_1};

endmodule




module ACS_col(clk,
			   rst,
			   data_id,
			   input_valid,
			   data_recv,
			   PM_in_1_1,
			   PM_in_1_2,
			   PM_in_2_1,
			   PM_in_2_2,
			   PM_in_3_1,
			   PM_in_3_2,
			   PM_in_4_1,
			   PM_in_4_2,
			   addr_in_1_1,
			   addr_in_1_2,
			   addr_in_2_1,
			   addr_in_2_2,
			   addr_in_3_1,
			   addr_in_3_2,
			   addr_in_4_1,
			   addr_in_4_2,
			   addr_out_1,
			   addr_out_2,
			   addr_out_3,
			   addr_out_4,
			   PM_out_1,
			   PM_out_2,
			   PM_out_3,
			   PM_out_4,
			   dec_out_1,
			   dec_out_2,
			   dec_out_3,
			   dec_out_4,
			   data_id_out,
			   data_rdy);
	
	input clk,rst,input_valid;
	input [1:0] data_recv,addr_in_1_1,addr_in_1_2,addr_in_2_1,addr_in_2_2,addr_in_3_1,addr_in_3_2,addr_in_4_1,addr_in_4_2;
	input [2:0] data_id;
	input [6:0] PM_in_1_1,PM_in_1_2,PM_in_2_1,PM_in_2_2,PM_in_3_1,PM_in_3_2,PM_in_4_1,PM_in_4_2;

	output dec_out_1,dec_out_2,dec_out_3,dec_out_4,data_rdy;
	output [1:0] addr_out_1,addr_out_2,addr_out_3,addr_out_4;
	output [2:0] data_id_out;
	output [6:0] PM_out_1,PM_out_2,PM_out_3,PM_out_4;

	//reg[1:0] self_state_1,self_state_2,self_state_3,self_state_4;

	//always begin
	//	self_state_1 = 2'b00;
	//	self_state_2 = 2'b01;
	//	self_state_3 = 2'b10;
	//	self_state_4 = 2'b11;
	//end

	ACS_module u_ACS_module_1(.clk(clk),
				  .rst(rst),
				  .data_id(data_id),
				  .self_state(2'b00),
				  .PM_in_1(PM_in_1_1),
				  .PM_in_2(PM_in_1_2),
				  .addr_in_1(addr_in_1_1),
				  .addr_in_2(addr_in_1_2),
				  .input_valid(input_valid),
				  .data_recv(data_recv),
				  .addr_out(addr_out_1),
				  .PM_out(PM_out_1),
				  .data_rdy(data_rdy),
				  .dec_out(dec_out_1),
				  .data_id_out(data_id_out));
	
	ACS_module u_ACS_module_2(.clk(clk),
				  .rst(rst),
				  .data_id(data_id),
				  .self_state(2'b01),
				  .PM_in_1(PM_in_2_1),
				  .PM_in_2(PM_in_2_2),
				  .addr_in_1(addr_in_2_1),
				  .addr_in_2(addr_in_2_2),
				  .input_valid(input_valid),
				  .data_recv(data_recv),
				  .addr_out(addr_out_2),
				  .PM_out(PM_out_2),
				  .data_rdy(data_rdy),
				  .dec_out(dec_out_2),
				  .data_id_out(data_id_out));
	
	ACS_module u_ACS_module_3(.clk(clk),
				  .rst(rst),
				  .data_id(data_id),
				  .self_state(2'b10),
				  .PM_in_1(PM_in_3_1),
				  .PM_in_2(PM_in_3_2),
				  .addr_in_1(addr_in_3_1),
				  .addr_in_2(addr_in_3_2),
				  .input_valid(input_valid),
				  .data_recv(data_recv),
				  .addr_out(addr_out_3),
				  .PM_out(PM_out_3),
				  .data_rdy(data_rdy),
				  .dec_out(dec_out_3),
				  .data_id_out(data_id_out));
	
	ACS_module u_ACS_module_4(.clk(clk),
				  .rst(rst),
				  .data_id(data_id),
				  .self_state(2'b11),
				  .PM_in_1(PM_in_4_1),
				  .PM_in_2(PM_in_4_2),
				  .addr_in_1(addr_in_4_1),
				  .addr_in_2(addr_in_4_2),
				  .input_valid(input_valid),
				  .data_recv(data_recv),
				  .addr_out(addr_out_4),
				  .PM_out(PM_out_4),
				  .data_rdy(data_rdy),
				  .dec_out(dec_out_4),
				  .data_id_out(data_id_out));

endmodule

// DONE BELOW

module ACS_module(clk,
				  rst,
				  data_id,
				  self_state,
				  PM_in_1,
				  term_1,
				  PM_in_2,
				  term_2,
				  addr_in_1,
				  addr_in_2,
				//  input_valid,
				  data_recv,
				  addr_out,
				  PM_out,
				  term_out,
				//  data_rdy,
				  dec_out,
				  data_id_out);

	input clk,rst,term_1,term_2;
	input [1:0] self_state,data_recv,addr_in_1,addr_in_2;
	input [2:0] data_id;
	input [6:0] PM_in_1,PM_in_2;

	output dec_out,term_out;
	output [1:0] addr_out;
	output [2:0] data_id_out;
	output [6:0] PM_out;

	wire w_term;
	wire [1:0] w_addr_out;
	wire [6:0] w_PM_out;



	ACS u_ACS(.self_state(self_state),
//		   .input_sig(input_valid),
		   .data_recv(data_recv),
		   .addr_in_1(addr_in_1),
		   .addr_in_2(addr_in_2),
		   .PMin1(PM_in_1),
		   .term_1(term_1),
		   .PMin2(PM_in_2),
		   .term_2(term_2),
		   .PMout(w_PM_out),
		   .term_out(w_term),
		   .addr_out(w_addr_out),
//		   .data_rdy(w_data_rdy),
		   .dec_out(w_dec_out));

	PM_mem u_PM_mem(.data_id(data_id),
			  .PM_clk(clk),
			  .PM_rst(rst),
		      .PM_in(w_PM_out),
		      .term_in(w_term),
//		      .data_en(w_data_rdy),
		      .addr_in(w_addr_out),
		      .dec_in(w_dec_out),
		      .PM_out(PM_out),
		      .term_out(term_out),
		      .addr_out(addr_out),
//		      .data_rdy(data_rdy),
		      .dec_out(dec_out),
		      .data_id_out(data_id_out));

endmodule