module ACS_matrix(clk,
				  rst,
				  data_recv_1,
				  data_recv_2,
				  data_recv_3,
				  data_recv_4,
				  data_recv_5,
				  data_recv_6,
				  data_recv_7,
				  data_recv_8,
				  data_out_1,
				  data_out_2,
				  data_out_3,
				  data_out_4,
				  PM_out_1,
				  PM_out_2,
				  PM_out_3,
				  PM_out_4);

	input clk,rst;
	input [1:0] data_recv_1,data_recv_2,data_recv_3,data_recv_4,data_recv_5,data_recv_6,data_recv_7,data_recv_8;

	output [6:0] PM_out_1,PM_out_2,PM_out_3,PM_out_4;
	output [7:0] data_out_1,data_out_2,data_out_3,data_out_4;

	wire [6:0] w_PM_1_to_2_1,w_PM_1_to_2_2,w_PM_1_to_2_3,w_PM_1_to_2_4,
			   w_PM_2_to_3_1,w_PM_2_to_3_2,w_PM_2_to_3_3,w_PM_2_to_3_4,
			   w_PM_3_to_4_1,w_PM_3_to_4_2,w_PM_3_to_4_3,w_PM_3_to_4_4,
			   w_PM_4_to_5_1,w_PM_4_to_5_2,w_PM_4_to_5_3,w_PM_4_to_5_4,
			   w_PM_5_to_6_1,w_PM_5_to_6_2,w_PM_5_to_6_3,w_PM_5_to_6_4,
			   w_PM_6_to_7_1,w_PM_6_to_7_2,w_PM_6_to_7_3,w_PM_6_to_7_4,
			   w_PM_7_to_8_1,w_PM_7_to_8_2,w_PM_7_to_8_3,w_PM_7_to_8_4;

	wire [7:0] w_data_1_to_2_1,w_data_1_to_2_2,w_data_1_to_2_3,w_data_1_to_2_4,
			   w_data_2_to_3_1,w_data_2_to_3_2,w_data_2_to_3_3,w_data_2_to_3_4,
			   w_data_3_to_4_1,w_data_3_to_4_2,w_data_3_to_4_3,w_data_3_to_4_4,
			   w_data_4_to_5_1,w_data_4_to_5_2,w_data_4_to_5_3,w_data_4_to_5_4,
			   w_data_5_to_6_1,w_data_5_to_6_2,w_data_5_to_6_3,w_data_5_to_6_4,
			   w_data_6_to_7_1,w_data_6_to_7_2,w_data_6_to_7_3,w_data_6_to_7_4,
			   w_data_7_to_8_1,w_data_7_to_8_2,w_data_7_to_8_3,w_data_7_to_8_4;

	ACS_col u_ACS_col_1(.clk(clk),
			   			.rst(rst),
			   			.data_recv(data_recv_1),
			   			.PM_in_1_1(7'b0),
			   			.PM_in_1_2(7'b0),
			   			.PM_in_2_1(7'b0),
			   			.PM_in_2_2(7'b0),
			   			.PM_in_3_1(7'b0),
			   			.PM_in_3_2(7'b0),
			   			.PM_in_4_1(7'b0),
			   			.PM_in_4_2(7'b0),
			   			.data_in_1_1(8'b0),
			   			.data_in_1_2(8'b0),
			   			.data_in_2_1(8'b0),
			   			.data_in_2_2(8'b0),
			   			.data_in_3_1(8'b0),
			   			.data_in_3_2(8'b0),
			   			.data_in_4_1(8'b0),
			   			.data_in_4_2(8'b0),
			   			.PM_out_1(w_PM_1_to_2_1),
			   			.PM_out_2(w_PM_1_to_2_2),
			   			.PM_out_3(w_PM_1_to_2_3),
			   			.PM_out_4(w_PM_1_to_2_4),
			   			.data_out_1(w_data_1_to_2_1),
			   			.data_out_2(w_data_1_to_2_2),
			   			.data_out_3(w_data_1_to_2_3),
		  				.data_out_4(w_data_1_to_2_4));

	ACS_col u_ACS_col_2(.clk(clk),
			   			.rst(rst),
			   			.data_recv(data_recv_2),
			   			.PM_in_1_1(w_PM_1_to_2_1),
			   			.PM_in_1_2(w_PM_1_to_2_2),
			   			.PM_in_2_1(w_PM_1_to_2_3),
			   			.PM_in_2_2(w_PM_1_to_2_4),
			   			.PM_in_3_1(w_PM_1_to_2_1),
			   			.PM_in_3_2(w_PM_1_to_2_2),
			   			.PM_in_4_1(w_PM_1_to_2_3),
			   			.PM_in_4_2(w_PM_1_to_2_4),
			   			.data_in_1_1(w_data_1_to_2_1),
			   			.data_in_1_2(w_data_1_to_2_2),
			   			.data_in_2_1(w_data_1_to_2_3),
			   			.data_in_2_2(w_data_1_to_2_4),
			   			.data_in_3_1(w_data_1_to_2_1),
			   			.data_in_3_2(w_data_1_to_2_2),
			   			.data_in_4_1(w_data_1_to_2_3),
			   			.data_in_4_2(w_data_1_to_2_4),
			   			.PM_out_1(w_PM_2_to_3_1),
			   			.PM_out_2(w_PM_2_to_3_2),
			   			.PM_out_3(w_PM_2_to_3_3),
			   			.PM_out_4(w_PM_2_to_3_4),
			   			.data_out_1(w_data_2_to_3_1),
			   			.data_out_2(w_data_2_to_3_2),
			   			.data_out_3(w_data_2_to_3_3),
		  				.data_out_4(w_data_2_to_3_4));

	ACS_col u_ACS_col_3(.clk(clk),
			   			.rst(rst),
			   			.data_recv(data_recv_3),
			   			.PM_in_1_1(w_PM_2_to_3_1),
			   			.PM_in_1_2(w_PM_2_to_3_2),
			   			.PM_in_2_1(w_PM_2_to_3_3),
			   			.PM_in_2_2(w_PM_2_to_3_4),
			   			.PM_in_3_1(w_PM_2_to_3_1),
			   			.PM_in_3_2(w_PM_2_to_3_2),
			   			.PM_in_4_1(w_PM_2_to_3_3),
			   			.PM_in_4_2(w_PM_2_to_3_4),
			   			.data_in_1_1(w_data_2_to_3_1),
			   			.data_in_1_2(w_data_2_to_3_2),
			   			.data_in_2_1(w_data_2_to_3_3),
			   			.data_in_2_2(w_data_2_to_3_4),
			   			.data_in_3_1(w_data_2_to_3_1),
			   			.data_in_3_2(w_data_2_to_3_2),
			   			.data_in_4_1(w_data_2_to_3_3),
			   			.data_in_4_2(w_data_2_to_3_4),
			   			.PM_out_1(w_PM_3_to_4_1),
			   			.PM_out_2(w_PM_3_to_4_2),
			   			.PM_out_3(w_PM_3_to_4_3),
			   			.PM_out_4(w_PM_3_to_4_4),
			   			.data_out_1(w_data_3_to_4_1),
			   			.data_out_2(w_data_3_to_4_2),
			   			.data_out_3(w_data_3_to_4_3),
		  				.data_out_4(w_data_3_to_4_4));

	ACS_col u_ACS_col_4(.clk(clk),
			   			.rst(rst),
			   			.data_recv(data_recv_4),
			   			.PM_in_1_1(w_PM_3_to_4_1),
			   			.PM_in_1_2(w_PM_3_to_4_2),
			   			.PM_in_2_1(w_PM_3_to_4_3),
			   			.PM_in_2_2(w_PM_3_to_4_4),
			   			.PM_in_3_1(w_PM_3_to_4_1),
			   			.PM_in_3_2(w_PM_3_to_4_2),
			   			.PM_in_4_1(w_PM_3_to_4_3),
			   			.PM_in_4_2(w_PM_3_to_4_4),
			   			.data_in_1_1(w_data_3_to_4_1),
			   			.data_in_1_2(w_data_3_to_4_2),
			   			.data_in_2_1(w_data_3_to_4_3),
			   			.data_in_2_2(w_data_3_to_4_4),
			   			.data_in_3_1(w_data_3_to_4_1),
			   			.data_in_3_2(w_data_3_to_4_2),
			   			.data_in_4_1(w_data_3_to_4_3),
			   			.data_in_4_2(w_data_3_to_4_4),
			   			.PM_out_1(w_PM_4_to_5_1),
			   			.PM_out_2(w_PM_4_to_5_2),
			   			.PM_out_3(w_PM_4_to_5_3),
			   			.PM_out_4(w_PM_4_to_5_4),
			   			.data_out_1(w_data_4_to_5_1),
			   			.data_out_2(w_data_4_to_5_2),
			   			.data_out_3(w_data_4_to_5_3),
		  				.data_out_4(w_data_4_to_5_4));

	ACS_col u_ACS_col_5(.clk(clk),
			   			.rst(rst),
			   			.data_recv(data_recv_5),
			   			.PM_in_1_1(w_PM_4_to_5_1),
			   			.PM_in_1_2(w_PM_4_to_5_2),
			   			.PM_in_2_1(w_PM_4_to_5_3),
			   			.PM_in_2_2(w_PM_4_to_5_4),
			   			.PM_in_3_1(w_PM_4_to_5_1),
			   			.PM_in_3_2(w_PM_4_to_5_2),
			   			.PM_in_4_1(w_PM_4_to_5_3),
			   			.PM_in_4_2(w_PM_4_to_5_4),
			   			.data_in_1_1(w_data_4_to_5_1),
			   			.data_in_1_2(w_data_4_to_5_2),
			   			.data_in_2_1(w_data_4_to_5_3),
			   			.data_in_2_2(w_data_4_to_5_4),
			   			.data_in_3_1(w_data_4_to_5_1),
			   			.data_in_3_2(w_data_4_to_5_2),
			   			.data_in_4_1(w_data_4_to_5_3),
			   			.data_in_4_2(w_data_4_to_5_4),
			   			.PM_out_1(w_PM_5_to_6_1),
			   			.PM_out_2(w_PM_5_to_6_2),
			   			.PM_out_3(w_PM_5_to_6_3),
			   			.PM_out_4(w_PM_5_to_6_4),
			   			.data_out_1(w_data_5_to_6_1),
			   			.data_out_2(w_data_5_to_6_2),
			   			.data_out_3(w_data_5_to_6_3),
		  				.data_out_4(w_data_5_to_6_4));

	ACS_col u_ACS_col_6(.clk(clk),
			   			.rst(rst),
			   			.data_recv(data_recv_6),
			   			.PM_in_1_1(w_PM_5_to_6_1),
			   			.PM_in_1_2(w_PM_5_to_6_2),
			   			.PM_in_2_1(w_PM_5_to_6_3),
			   			.PM_in_2_2(w_PM_5_to_6_4),
			   			.PM_in_3_1(w_PM_5_to_6_1),
			   			.PM_in_3_2(w_PM_5_to_6_2),
			   			.PM_in_4_1(w_PM_5_to_6_3),
			   			.PM_in_4_2(w_PM_5_to_6_4),
			   			.data_in_1_1(w_data_5_to_6_1),
			   			.data_in_1_2(w_data_5_to_6_2),
			   			.data_in_2_1(w_data_5_to_6_3),
			   			.data_in_2_2(w_data_5_to_6_4),
			   			.data_in_3_1(w_data_5_to_6_1),
			   			.data_in_3_2(w_data_5_to_6_2),
			   			.data_in_4_1(w_data_5_to_6_3),
			   			.data_in_4_2(w_data_5_to_6_4),
			   			.PM_out_1(w_PM_6_to_7_1),
			   			.PM_out_2(w_PM_6_to_7_2),
			   			.PM_out_3(w_PM_6_to_7_3),
			   			.PM_out_4(w_PM_6_to_7_4),
			   			.data_out_1(w_data_6_to_7_1),
			   			.data_out_2(w_data_6_to_7_2),
			   			.data_out_3(w_data_6_to_7_3),
		  				.data_out_4(w_data_6_to_7_4));

	ACS_col u_ACS_col_7(.clk(clk),
			   			.rst(rst),
			   			.data_recv(data_recv_7),
			   			.PM_in_1_1(w_PM_6_to_7_1),
			   			.PM_in_1_2(w_PM_6_to_7_2),
			   			.PM_in_2_1(w_PM_6_to_7_3),
			   			.PM_in_2_2(w_PM_6_to_7_4),
			   			.PM_in_3_1(w_PM_6_to_7_1),
			   			.PM_in_3_2(w_PM_6_to_7_2),
			   			.PM_in_4_1(w_PM_6_to_7_3),
			   			.PM_in_4_2(w_PM_6_to_7_4),
			   			.data_in_1_1(w_data_6_to_7_1),
			   			.data_in_1_2(w_data_6_to_7_2),
			   			.data_in_2_1(w_data_6_to_7_3),
			   			.data_in_2_2(w_data_6_to_7_4),
			   			.data_in_3_1(w_data_6_to_7_1),
			   			.data_in_3_2(w_data_6_to_7_2),
			   			.data_in_4_1(w_data_6_to_7_3),
			   			.data_in_4_2(w_data_6_to_7_4),
			   			.PM_out_1(w_PM_7_to_8_1),
			   			.PM_out_2(w_PM_7_to_8_2),
			   			.PM_out_3(w_PM_7_to_8_3),
			   			.PM_out_4(w_PM_7_to_8_4),
			   			.data_out_1(w_data_7_to_8_1),
			   			.data_out_2(w_data_7_to_8_2),
			   			.data_out_3(w_data_7_to_8_3),
		  				.data_out_4(w_data_7_to_8_4));

	ACS_col u_ACS_col_8(.clk(clk),
			   			.rst(rst),
			   			.data_recv(data_recv_8),
			   			.PM_in_1_1(w_PM_7_to_8_1),
			   			.PM_in_1_2(w_PM_7_to_8_2),
			   			.PM_in_2_1(w_PM_7_to_8_3),
			   			.PM_in_2_2(w_PM_7_to_8_4),
			   			.PM_in_3_1(w_PM_7_to_8_1),
			   			.PM_in_3_2(w_PM_7_to_8_2),
			   			.PM_in_4_1(w_PM_7_to_8_3),
			   			.PM_in_4_2(w_PM_7_to_8_4),
			   			.data_in_1_1(w_data_7_to_8_1),
			   			.data_in_1_2(w_data_7_to_8_2),
			   			.data_in_2_1(w_data_7_to_8_3),
			   			.data_in_2_2(w_data_7_to_8_4),
			   			.data_in_3_1(w_data_7_to_8_1),
			   			.data_in_3_2(w_data_7_to_8_2),
			   			.data_in_4_1(w_data_7_to_8_3),
			   			.data_in_4_2(w_data_7_to_8_4),
			   			.PM_out_1(PM_out_1),
			   			.PM_out_2(PM_out_2),
			   			.PM_out_3(PM_out_3),
			   			.PM_out_4(PM_out_4),
			   			.data_out_1(data_out_1),
			   			.data_out_2(data_out_2),
			   			.data_out_3(data_out_3),
		  				.data_out_4(data_out_4));

endmodule

module ACS_col(clk,
			   rst,
			   data_recv,
			   PM_in_1_1,
			   PM_in_1_2,
			   PM_in_2_1,
			   PM_in_2_2,
			   PM_in_3_1,
			   PM_in_3_2,
			   PM_in_4_1,
			   PM_in_4_2,
			   data_in_1_1,
			   data_in_1_2,
			   data_in_2_1,
			   data_in_2_2,
			   data_in_3_1,
			   data_in_3_2,
			   data_in_4_1,
			   data_in_4_2,
			   PM_out_1,
			   PM_out_2,
			   PM_out_3,
			   PM_out_4,
			   data_out_1,
			   data_out_2,
			   data_out_3,
			   data_out_4);
	
	input clk,rst;
	input [1:0] data_recv;
	input [6:0] PM_in_1_1,PM_in_1_2,PM_in_2_1,PM_in_2_2,PM_in_3_1,PM_in_3_2,PM_in_4_1,PM_in_4_2;
	input [7:0] data_in_1_1,data_in_1_2,data_in_2_1,data_in_2_2,data_in_3_1,data_in_3_2,data_in_4_1,data_in_4_2;

	output [6:0] PM_out_1,PM_out_2,PM_out_3,PM_out_4;
	output [7:0] data_out_1,data_out_2,data_out_3,data_out_4;

	//module ACS_mem(rst,
	//		   clk,
	//		   self_state,
	//		   data_recv,
	//		   PM_in_1,
	//		   PM_in_2,
	//		   data_in_1,
	//		   data_in_2,
	//		   PM_out,
	//		   data_out);

	ACS_mem u_ACS_mem_1(.rst(rst),
						.clk(clk),
				 		.self_state(2'b00),
				 		.data_recv(data_recv),
				  		.PM_in_1(PM_in_1_1),
				  		.PM_in_2(PM_in_1_2),
				  		.data_in_1(data_in_1_1),
				  		.data_in_2(data_in_1_2),
				  		.PM_out(PM_out_1),
				  		.data_out(data_out_1));

	ACS_mem u_ACS_mem_2(.rst(rst),
						.clk(clk),
				 		.self_state(2'b01),
				 		.data_recv(data_recv),
				  		.PM_in_1(PM_in_2_1),
				  		.PM_in_2(PM_in_2_2),
				  		.data_in_1(data_in_2_1),
				  		.data_in_2(data_in_2_2),
				  		.PM_out(PM_out_2),
				  		.data_out(data_out_2));

	ACS_mem u_ACS_mem_3(.rst(rst),
						.clk(clk),
				 		.self_state(2'b10),
				 		.data_recv(data_recv),
				  		.PM_in_1(PM_in_3_1),
				  		.PM_in_2(PM_in_3_2),
				  		.data_in_1(data_in_3_1),
				  		.data_in_2(data_in_3_2),
				  		.PM_out(PM_out_3),
				  		.data_out(data_out_3));

	ACS_mem u_ACS_mem_4(.rst(rst),
						.clk(clk),
				 		.self_state(2'b11),
				 		.data_recv(data_recv),
				  		.PM_in_1(PM_in_4_1),
				  		.PM_in_2(PM_in_4_2),
				  		.data_in_1(data_in_4_1),
				  		.data_in_2(data_in_4_2),
				  		.PM_out(PM_out_4),
				  		.data_out(data_out_4));

endmodule